netcdf var4d {
dimensions:
	time = 3 ;
	level = 2 ;
	lat = 4 ;
	lon = 5 ;
variables:
	float temp_surface(lat, lon) ;
	float temp_profile(time, lat, lon) ;
	float temp_3d(time, level, lat, lon) ;
data:

 temp_surface =
  273.15, 275.15, 277.15, 279.15, 281.15,
  278.15, 280.15, 282.15, 284.15, 286.15,
  283.15, 285.15, 287.15, 289.15, 291.15,
  288.15, 290.15, 292.15, 294.15, 296.15 ;

 temp_profile =
  273.15, 275.15, 277.15, 279.15, 281.15,
  278.15, 280.15, 282.15, 284.15, 286.15,
  283.15, 285.15, 287.15, 289.15, 291.15,
  288.15, 290.15, 292.15, 294.15, 296.15,
  274.15, 276.15, 278.15, 280.15, 282.15,
  279.15, 281.15, 283.15, 285.15, 287.15,
  284.15, 286.15, 288.15, 290.15, 292.15,
  289.15, 291.15, 293.15, 295.15, 297.15,
  275.15, 277.15, 279.15, 281.15, 283.15,
  280.15, 282.15, 284.15, 286.15, 288.15,
  285.15, 287.15, 289.15, 291.15, 293.15,
  290.15, 292.15, 294.15, 296.15, 298.15 ;

 temp_3d =
  273.15, 275.15, 277.15, 279.15, 281.15,
  278.15, 280.15, 282.15, 284.15, 286.15,
  283.15, 285.15, 287.15, 289.15, 291.15,
  288.15, 290.15, 292.15, 294.15, 296.15,
  283.15, 285.15, 287.15, 289.15, 291.15,
  288.15, 290.15, 292.15, 294.15, 296.15,
  293.15, 295.15, 297.15, 299.15, 301.15,
  298.15, 300.15, 302.15, 304.15, 306.15,
  274.15, 276.15, 278.15, 280.15, 282.15,
  279.15, 281.15, 283.15, 285.15, 287.15,
  284.15, 286.15, 288.15, 290.15, 292.15,
  289.15, 291.15, 293.15, 295.15, 297.15,
  284.15, 286.15, 288.15, 290.15, 292.15,
  289.15, 291.15, 293.15, 295.15, 297.15,
  294.15, 296.15, 298.15, 300.15, 302.15,
  299.15, 301.15, 303.15, 305.15, 307.15,
  275.15, 277.15, 279.15, 281.15, 283.15,
  280.15, 282.15, 284.15, 286.15, 288.15,
  285.15, 287.15, 289.15, 291.15, 293.15,
  290.15, 292.15, 294.15, 296.15, 298.15,
  285.15, 287.15, 289.15, 291.15, 293.15,
  290.15, 292.15, 294.15, 296.15, 298.15,
  295.15, 297.15, 299.15, 301.15, 303.15,
  300.15, 302.15, 304.15, 306.15, 308.15 ;
}
