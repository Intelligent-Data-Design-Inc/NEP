netcdf format_netcdf4 {
dimensions:
	time = 10 ;
	lat = 20 ;
	lon = 30 ;
variables:
	float temperature(time, lat, lon) ;
		temperature:units = "K" ;
	float pressure(time, lat, lon) ;
		pressure:units = "hPa" ;
data:

 temperature =
  273.15, 273.35, 273.55, 273.75, 273.95, 274.15, 274.35, 274.55, 274.75, 
    274.95, 275.15, 275.35, 275.55, 275.75, 275.95, 276.15, 276.35, 276.55, 
    276.75, 276.95, 277.15, 277.35, 277.55, 277.75, 277.95, 278.15, 278.35, 
    278.55, 278.75, 278.95,
  273.65, 273.85, 274.05, 274.25, 274.45, 274.65, 274.85, 275.05, 275.25, 
    275.45, 275.65, 275.85, 276.05, 276.25, 276.45, 276.65, 276.85, 277.05, 
    277.25, 277.45, 277.65, 277.85, 278.05, 278.25, 278.45, 278.65, 278.85, 
    279.05, 279.25, 279.45,
  274.15, 274.35, 274.55, 274.75, 274.95, 275.15, 275.35, 275.55, 275.75, 
    275.95, 276.15, 276.35, 276.55, 276.75, 276.95, 277.15, 277.35, 277.55, 
    277.75, 277.95, 278.15, 278.35, 278.55, 278.75, 278.95, 279.15, 279.35, 
    279.55, 279.75, 279.95,
  274.65, 274.85, 275.05, 275.25, 275.45, 275.65, 275.85, 276.05, 276.25, 
    276.45, 276.65, 276.85, 277.05, 277.25, 277.45, 277.65, 277.85, 278.05, 
    278.25, 278.45, 278.65, 278.85, 279.05, 279.25, 279.45, 279.65, 279.85, 
    280.05, 280.25, 280.45,
  275.15, 275.35, 275.55, 275.75, 275.95, 276.15, 276.35, 276.55, 276.75, 
    276.95, 277.15, 277.35, 277.55, 277.75, 277.95, 278.15, 278.35, 278.55, 
    278.75, 278.95, 279.15, 279.35, 279.55, 279.75, 279.95, 280.15, 280.35, 
    280.55, 280.75, 280.95,
  275.65, 275.85, 276.05, 276.25, 276.45, 276.65, 276.85, 277.05, 277.25, 
    277.45, 277.65, 277.85, 278.05, 278.25, 278.45, 278.65, 278.85, 279.05, 
    279.25, 279.45, 279.65, 279.85, 280.05, 280.25, 280.45, 280.65, 280.85, 
    281.05, 281.25, 281.45,
  276.15, 276.35, 276.55, 276.75, 276.95, 277.15, 277.35, 277.55, 277.75, 
    277.95, 278.15, 278.35, 278.55, 278.75, 278.95, 279.15, 279.35, 279.55, 
    279.75, 279.95, 280.15, 280.35, 280.55, 280.75, 280.95, 281.15, 281.35, 
    281.55, 281.75, 281.95,
  276.65, 276.85, 277.05, 277.25, 277.45, 277.65, 277.85, 278.05, 278.25, 
    278.45, 278.65, 278.85, 279.05, 279.25, 279.45, 279.65, 279.85, 280.05, 
    280.25, 280.45, 280.65, 280.85, 281.05, 281.25, 281.45, 281.65, 281.85, 
    282.05, 282.25, 282.45,
  277.15, 277.35, 277.55, 277.75, 277.95, 278.15, 278.35, 278.55, 278.75, 
    278.95, 279.15, 279.35, 279.55, 279.75, 279.95, 280.15, 280.35, 280.55, 
    280.75, 280.95, 281.15, 281.35, 281.55, 281.75, 281.95, 282.15, 282.35, 
    282.55, 282.75, 282.95,
  277.65, 277.85, 278.05, 278.25, 278.45, 278.65, 278.85, 279.05, 279.25, 
    279.45, 279.65, 279.85, 280.05, 280.25, 280.45, 280.65, 280.85, 281.05, 
    281.25, 281.45, 281.65, 281.85, 282.05, 282.25, 282.45, 282.65, 282.85, 
    283.05, 283.25, 283.45,
  278.15, 278.35, 278.55, 278.75, 278.95, 279.15, 279.35, 279.55, 279.75, 
    279.95, 280.15, 280.35, 280.55, 280.75, 280.95, 281.15, 281.35, 281.55, 
    281.75, 281.95, 282.15, 282.35, 282.55, 282.75, 282.95, 283.15, 283.35, 
    283.55, 283.75, 283.95,
  278.65, 278.85, 279.05, 279.25, 279.45, 279.65, 279.85, 280.05, 280.25, 
    280.45, 280.65, 280.85, 281.05, 281.25, 281.45, 281.65, 281.85, 282.05, 
    282.25, 282.45, 282.65, 282.85, 283.05, 283.25, 283.45, 283.65, 283.85, 
    284.05, 284.25, 284.45,
  279.15, 279.35, 279.55, 279.75, 279.95, 280.15, 280.35, 280.55, 280.75, 
    280.95, 281.15, 281.35, 281.55, 281.75, 281.95, 282.15, 282.35, 282.55, 
    282.75, 282.95, 283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 
    284.55, 284.75, 284.95,
  279.65, 279.85, 280.05, 280.25, 280.45, 280.65, 280.85, 281.05, 281.25, 
    281.45, 281.65, 281.85, 282.05, 282.25, 282.45, 282.65, 282.85, 283.05, 
    283.25, 283.45, 283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 
    285.05, 285.25, 285.45,
  280.15, 280.35, 280.55, 280.75, 280.95, 281.15, 281.35, 281.55, 281.75, 
    281.95, 282.15, 282.35, 282.55, 282.75, 282.95, 283.15, 283.35, 283.55, 
    283.75, 283.95, 284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 
    285.55, 285.75, 285.95,
  280.65, 280.85, 281.05, 281.25, 281.45, 281.65, 281.85, 282.05, 282.25, 
    282.45, 282.65, 282.85, 283.05, 283.25, 283.45, 283.65, 283.85, 284.05, 
    284.25, 284.45, 284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 
    286.05, 286.25, 286.45,
  281.15, 281.35, 281.55, 281.75, 281.95, 282.15, 282.35, 282.55, 282.75, 
    282.95, 283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 284.55, 
    284.75, 284.95, 285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 
    286.55, 286.75, 286.95,
  281.65, 281.85, 282.05, 282.25, 282.45, 282.65, 282.85, 283.05, 283.25, 
    283.45, 283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 285.05, 
    285.25, 285.45, 285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 
    287.05, 287.25, 287.45,
  282.15, 282.35, 282.55, 282.75, 282.95, 283.15, 283.35, 283.55, 283.75, 
    283.95, 284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 285.55, 
    285.75, 285.95, 286.15, 286.35, 286.55, 286.75, 286.95, 287.15, 287.35, 
    287.55, 287.75, 287.95,
  282.65, 282.85, 283.05, 283.25, 283.45, 283.65, 283.85, 284.05, 284.25, 
    284.45, 284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 286.05, 
    286.25, 286.45, 286.65, 286.85, 287.05, 287.25, 287.45, 287.65, 287.85, 
    288.05, 288.25, 288.45,
  274.15, 274.35, 274.55, 274.75, 274.95, 275.15, 275.35, 275.55, 275.75, 
    275.95, 276.15, 276.35, 276.55, 276.75, 276.95, 277.15, 277.35, 277.55, 
    277.75, 277.95, 278.15, 278.35, 278.55, 278.75, 278.95, 279.15, 279.35, 
    279.55, 279.75, 279.95,
  274.65, 274.85, 275.05, 275.25, 275.45, 275.65, 275.85, 276.05, 276.25, 
    276.45, 276.65, 276.85, 277.05, 277.25, 277.45, 277.65, 277.85, 278.05, 
    278.25, 278.45, 278.65, 278.85, 279.05, 279.25, 279.45, 279.65, 279.85, 
    280.05, 280.25, 280.45,
  275.15, 275.35, 275.55, 275.75, 275.95, 276.15, 276.35, 276.55, 276.75, 
    276.95, 277.15, 277.35, 277.55, 277.75, 277.95, 278.15, 278.35, 278.55, 
    278.75, 278.95, 279.15, 279.35, 279.55, 279.75, 279.95, 280.15, 280.35, 
    280.55, 280.75, 280.95,
  275.65, 275.85, 276.05, 276.25, 276.45, 276.65, 276.85, 277.05, 277.25, 
    277.45, 277.65, 277.85, 278.05, 278.25, 278.45, 278.65, 278.85, 279.05, 
    279.25, 279.45, 279.65, 279.85, 280.05, 280.25, 280.45, 280.65, 280.85, 
    281.05, 281.25, 281.45,
  276.15, 276.35, 276.55, 276.75, 276.95, 277.15, 277.35, 277.55, 277.75, 
    277.95, 278.15, 278.35, 278.55, 278.75, 278.95, 279.15, 279.35, 279.55, 
    279.75, 279.95, 280.15, 280.35, 280.55, 280.75, 280.95, 281.15, 281.35, 
    281.55, 281.75, 281.95,
  276.65, 276.85, 277.05, 277.25, 277.45, 277.65, 277.85, 278.05, 278.25, 
    278.45, 278.65, 278.85, 279.05, 279.25, 279.45, 279.65, 279.85, 280.05, 
    280.25, 280.45, 280.65, 280.85, 281.05, 281.25, 281.45, 281.65, 281.85, 
    282.05, 282.25, 282.45,
  277.15, 277.35, 277.55, 277.75, 277.95, 278.15, 278.35, 278.55, 278.75, 
    278.95, 279.15, 279.35, 279.55, 279.75, 279.95, 280.15, 280.35, 280.55, 
    280.75, 280.95, 281.15, 281.35, 281.55, 281.75, 281.95, 282.15, 282.35, 
    282.55, 282.75, 282.95,
  277.65, 277.85, 278.05, 278.25, 278.45, 278.65, 278.85, 279.05, 279.25, 
    279.45, 279.65, 279.85, 280.05, 280.25, 280.45, 280.65, 280.85, 281.05, 
    281.25, 281.45, 281.65, 281.85, 282.05, 282.25, 282.45, 282.65, 282.85, 
    283.05, 283.25, 283.45,
  278.15, 278.35, 278.55, 278.75, 278.95, 279.15, 279.35, 279.55, 279.75, 
    279.95, 280.15, 280.35, 280.55, 280.75, 280.95, 281.15, 281.35, 281.55, 
    281.75, 281.95, 282.15, 282.35, 282.55, 282.75, 282.95, 283.15, 283.35, 
    283.55, 283.75, 283.95,
  278.65, 278.85, 279.05, 279.25, 279.45, 279.65, 279.85, 280.05, 280.25, 
    280.45, 280.65, 280.85, 281.05, 281.25, 281.45, 281.65, 281.85, 282.05, 
    282.25, 282.45, 282.65, 282.85, 283.05, 283.25, 283.45, 283.65, 283.85, 
    284.05, 284.25, 284.45,
  279.15, 279.35, 279.55, 279.75, 279.95, 280.15, 280.35, 280.55, 280.75, 
    280.95, 281.15, 281.35, 281.55, 281.75, 281.95, 282.15, 282.35, 282.55, 
    282.75, 282.95, 283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 
    284.55, 284.75, 284.95,
  279.65, 279.85, 280.05, 280.25, 280.45, 280.65, 280.85, 281.05, 281.25, 
    281.45, 281.65, 281.85, 282.05, 282.25, 282.45, 282.65, 282.85, 283.05, 
    283.25, 283.45, 283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 
    285.05, 285.25, 285.45,
  280.15, 280.35, 280.55, 280.75, 280.95, 281.15, 281.35, 281.55, 281.75, 
    281.95, 282.15, 282.35, 282.55, 282.75, 282.95, 283.15, 283.35, 283.55, 
    283.75, 283.95, 284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 
    285.55, 285.75, 285.95,
  280.65, 280.85, 281.05, 281.25, 281.45, 281.65, 281.85, 282.05, 282.25, 
    282.45, 282.65, 282.85, 283.05, 283.25, 283.45, 283.65, 283.85, 284.05, 
    284.25, 284.45, 284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 
    286.05, 286.25, 286.45,
  281.15, 281.35, 281.55, 281.75, 281.95, 282.15, 282.35, 282.55, 282.75, 
    282.95, 283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 284.55, 
    284.75, 284.95, 285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 
    286.55, 286.75, 286.95,
  281.65, 281.85, 282.05, 282.25, 282.45, 282.65, 282.85, 283.05, 283.25, 
    283.45, 283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 285.05, 
    285.25, 285.45, 285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 
    287.05, 287.25, 287.45,
  282.15, 282.35, 282.55, 282.75, 282.95, 283.15, 283.35, 283.55, 283.75, 
    283.95, 284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 285.55, 
    285.75, 285.95, 286.15, 286.35, 286.55, 286.75, 286.95, 287.15, 287.35, 
    287.55, 287.75, 287.95,
  282.65, 282.85, 283.05, 283.25, 283.45, 283.65, 283.85, 284.05, 284.25, 
    284.45, 284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 286.05, 
    286.25, 286.45, 286.65, 286.85, 287.05, 287.25, 287.45, 287.65, 287.85, 
    288.05, 288.25, 288.45,
  283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 284.55, 284.75, 
    284.95, 285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 286.55, 
    286.75, 286.95, 287.15, 287.35, 287.55, 287.75, 287.95, 288.15, 288.35, 
    288.55, 288.75, 288.95,
  283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 285.05, 285.25, 
    285.45, 285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 287.05, 
    287.25, 287.45, 287.65, 287.85, 288.05, 288.25, 288.45, 288.65, 288.85, 
    289.05, 289.25, 289.45,
  275.15, 275.35, 275.55, 275.75, 275.95, 276.15, 276.35, 276.55, 276.75, 
    276.95, 277.15, 277.35, 277.55, 277.75, 277.95, 278.15, 278.35, 278.55, 
    278.75, 278.95, 279.15, 279.35, 279.55, 279.75, 279.95, 280.15, 280.35, 
    280.55, 280.75, 280.95,
  275.65, 275.85, 276.05, 276.25, 276.45, 276.65, 276.85, 277.05, 277.25, 
    277.45, 277.65, 277.85, 278.05, 278.25, 278.45, 278.65, 278.85, 279.05, 
    279.25, 279.45, 279.65, 279.85, 280.05, 280.25, 280.45, 280.65, 280.85, 
    281.05, 281.25, 281.45,
  276.15, 276.35, 276.55, 276.75, 276.95, 277.15, 277.35, 277.55, 277.75, 
    277.95, 278.15, 278.35, 278.55, 278.75, 278.95, 279.15, 279.35, 279.55, 
    279.75, 279.95, 280.15, 280.35, 280.55, 280.75, 280.95, 281.15, 281.35, 
    281.55, 281.75, 281.95,
  276.65, 276.85, 277.05, 277.25, 277.45, 277.65, 277.85, 278.05, 278.25, 
    278.45, 278.65, 278.85, 279.05, 279.25, 279.45, 279.65, 279.85, 280.05, 
    280.25, 280.45, 280.65, 280.85, 281.05, 281.25, 281.45, 281.65, 281.85, 
    282.05, 282.25, 282.45,
  277.15, 277.35, 277.55, 277.75, 277.95, 278.15, 278.35, 278.55, 278.75, 
    278.95, 279.15, 279.35, 279.55, 279.75, 279.95, 280.15, 280.35, 280.55, 
    280.75, 280.95, 281.15, 281.35, 281.55, 281.75, 281.95, 282.15, 282.35, 
    282.55, 282.75, 282.95,
  277.65, 277.85, 278.05, 278.25, 278.45, 278.65, 278.85, 279.05, 279.25, 
    279.45, 279.65, 279.85, 280.05, 280.25, 280.45, 280.65, 280.85, 281.05, 
    281.25, 281.45, 281.65, 281.85, 282.05, 282.25, 282.45, 282.65, 282.85, 
    283.05, 283.25, 283.45,
  278.15, 278.35, 278.55, 278.75, 278.95, 279.15, 279.35, 279.55, 279.75, 
    279.95, 280.15, 280.35, 280.55, 280.75, 280.95, 281.15, 281.35, 281.55, 
    281.75, 281.95, 282.15, 282.35, 282.55, 282.75, 282.95, 283.15, 283.35, 
    283.55, 283.75, 283.95,
  278.65, 278.85, 279.05, 279.25, 279.45, 279.65, 279.85, 280.05, 280.25, 
    280.45, 280.65, 280.85, 281.05, 281.25, 281.45, 281.65, 281.85, 282.05, 
    282.25, 282.45, 282.65, 282.85, 283.05, 283.25, 283.45, 283.65, 283.85, 
    284.05, 284.25, 284.45,
  279.15, 279.35, 279.55, 279.75, 279.95, 280.15, 280.35, 280.55, 280.75, 
    280.95, 281.15, 281.35, 281.55, 281.75, 281.95, 282.15, 282.35, 282.55, 
    282.75, 282.95, 283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 
    284.55, 284.75, 284.95,
  279.65, 279.85, 280.05, 280.25, 280.45, 280.65, 280.85, 281.05, 281.25, 
    281.45, 281.65, 281.85, 282.05, 282.25, 282.45, 282.65, 282.85, 283.05, 
    283.25, 283.45, 283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 
    285.05, 285.25, 285.45,
  280.15, 280.35, 280.55, 280.75, 280.95, 281.15, 281.35, 281.55, 281.75, 
    281.95, 282.15, 282.35, 282.55, 282.75, 282.95, 283.15, 283.35, 283.55, 
    283.75, 283.95, 284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 
    285.55, 285.75, 285.95,
  280.65, 280.85, 281.05, 281.25, 281.45, 281.65, 281.85, 282.05, 282.25, 
    282.45, 282.65, 282.85, 283.05, 283.25, 283.45, 283.65, 283.85, 284.05, 
    284.25, 284.45, 284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 
    286.05, 286.25, 286.45,
  281.15, 281.35, 281.55, 281.75, 281.95, 282.15, 282.35, 282.55, 282.75, 
    282.95, 283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 284.55, 
    284.75, 284.95, 285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 
    286.55, 286.75, 286.95,
  281.65, 281.85, 282.05, 282.25, 282.45, 282.65, 282.85, 283.05, 283.25, 
    283.45, 283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 285.05, 
    285.25, 285.45, 285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 
    287.05, 287.25, 287.45,
  282.15, 282.35, 282.55, 282.75, 282.95, 283.15, 283.35, 283.55, 283.75, 
    283.95, 284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 285.55, 
    285.75, 285.95, 286.15, 286.35, 286.55, 286.75, 286.95, 287.15, 287.35, 
    287.55, 287.75, 287.95,
  282.65, 282.85, 283.05, 283.25, 283.45, 283.65, 283.85, 284.05, 284.25, 
    284.45, 284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 286.05, 
    286.25, 286.45, 286.65, 286.85, 287.05, 287.25, 287.45, 287.65, 287.85, 
    288.05, 288.25, 288.45,
  283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 284.55, 284.75, 
    284.95, 285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 286.55, 
    286.75, 286.95, 287.15, 287.35, 287.55, 287.75, 287.95, 288.15, 288.35, 
    288.55, 288.75, 288.95,
  283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 285.05, 285.25, 
    285.45, 285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 287.05, 
    287.25, 287.45, 287.65, 287.85, 288.05, 288.25, 288.45, 288.65, 288.85, 
    289.05, 289.25, 289.45,
  284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 285.55, 285.75, 
    285.95, 286.15, 286.35, 286.55, 286.75, 286.95, 287.15, 287.35, 287.55, 
    287.75, 287.95, 288.15, 288.35, 288.55, 288.75, 288.95, 289.15, 289.35, 
    289.55, 289.75, 289.95,
  284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 286.05, 286.25, 
    286.45, 286.65, 286.85, 287.05, 287.25, 287.45, 287.65, 287.85, 288.05, 
    288.25, 288.45, 288.65, 288.85, 289.05, 289.25, 289.45, 289.65, 289.85, 
    290.05, 290.25, 290.45,
  276.15, 276.35, 276.55, 276.75, 276.95, 277.15, 277.35, 277.55, 277.75, 
    277.95, 278.15, 278.35, 278.55, 278.75, 278.95, 279.15, 279.35, 279.55, 
    279.75, 279.95, 280.15, 280.35, 280.55, 280.75, 280.95, 281.15, 281.35, 
    281.55, 281.75, 281.95,
  276.65, 276.85, 277.05, 277.25, 277.45, 277.65, 277.85, 278.05, 278.25, 
    278.45, 278.65, 278.85, 279.05, 279.25, 279.45, 279.65, 279.85, 280.05, 
    280.25, 280.45, 280.65, 280.85, 281.05, 281.25, 281.45, 281.65, 281.85, 
    282.05, 282.25, 282.45,
  277.15, 277.35, 277.55, 277.75, 277.95, 278.15, 278.35, 278.55, 278.75, 
    278.95, 279.15, 279.35, 279.55, 279.75, 279.95, 280.15, 280.35, 280.55, 
    280.75, 280.95, 281.15, 281.35, 281.55, 281.75, 281.95, 282.15, 282.35, 
    282.55, 282.75, 282.95,
  277.65, 277.85, 278.05, 278.25, 278.45, 278.65, 278.85, 279.05, 279.25, 
    279.45, 279.65, 279.85, 280.05, 280.25, 280.45, 280.65, 280.85, 281.05, 
    281.25, 281.45, 281.65, 281.85, 282.05, 282.25, 282.45, 282.65, 282.85, 
    283.05, 283.25, 283.45,
  278.15, 278.35, 278.55, 278.75, 278.95, 279.15, 279.35, 279.55, 279.75, 
    279.95, 280.15, 280.35, 280.55, 280.75, 280.95, 281.15, 281.35, 281.55, 
    281.75, 281.95, 282.15, 282.35, 282.55, 282.75, 282.95, 283.15, 283.35, 
    283.55, 283.75, 283.95,
  278.65, 278.85, 279.05, 279.25, 279.45, 279.65, 279.85, 280.05, 280.25, 
    280.45, 280.65, 280.85, 281.05, 281.25, 281.45, 281.65, 281.85, 282.05, 
    282.25, 282.45, 282.65, 282.85, 283.05, 283.25, 283.45, 283.65, 283.85, 
    284.05, 284.25, 284.45,
  279.15, 279.35, 279.55, 279.75, 279.95, 280.15, 280.35, 280.55, 280.75, 
    280.95, 281.15, 281.35, 281.55, 281.75, 281.95, 282.15, 282.35, 282.55, 
    282.75, 282.95, 283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 
    284.55, 284.75, 284.95,
  279.65, 279.85, 280.05, 280.25, 280.45, 280.65, 280.85, 281.05, 281.25, 
    281.45, 281.65, 281.85, 282.05, 282.25, 282.45, 282.65, 282.85, 283.05, 
    283.25, 283.45, 283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 
    285.05, 285.25, 285.45,
  280.15, 280.35, 280.55, 280.75, 280.95, 281.15, 281.35, 281.55, 281.75, 
    281.95, 282.15, 282.35, 282.55, 282.75, 282.95, 283.15, 283.35, 283.55, 
    283.75, 283.95, 284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 
    285.55, 285.75, 285.95,
  280.65, 280.85, 281.05, 281.25, 281.45, 281.65, 281.85, 282.05, 282.25, 
    282.45, 282.65, 282.85, 283.05, 283.25, 283.45, 283.65, 283.85, 284.05, 
    284.25, 284.45, 284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 
    286.05, 286.25, 286.45,
  281.15, 281.35, 281.55, 281.75, 281.95, 282.15, 282.35, 282.55, 282.75, 
    282.95, 283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 284.55, 
    284.75, 284.95, 285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 
    286.55, 286.75, 286.95,
  281.65, 281.85, 282.05, 282.25, 282.45, 282.65, 282.85, 283.05, 283.25, 
    283.45, 283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 285.05, 
    285.25, 285.45, 285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 
    287.05, 287.25, 287.45,
  282.15, 282.35, 282.55, 282.75, 282.95, 283.15, 283.35, 283.55, 283.75, 
    283.95, 284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 285.55, 
    285.75, 285.95, 286.15, 286.35, 286.55, 286.75, 286.95, 287.15, 287.35, 
    287.55, 287.75, 287.95,
  282.65, 282.85, 283.05, 283.25, 283.45, 283.65, 283.85, 284.05, 284.25, 
    284.45, 284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 286.05, 
    286.25, 286.45, 286.65, 286.85, 287.05, 287.25, 287.45, 287.65, 287.85, 
    288.05, 288.25, 288.45,
  283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 284.55, 284.75, 
    284.95, 285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 286.55, 
    286.75, 286.95, 287.15, 287.35, 287.55, 287.75, 287.95, 288.15, 288.35, 
    288.55, 288.75, 288.95,
  283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 285.05, 285.25, 
    285.45, 285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 287.05, 
    287.25, 287.45, 287.65, 287.85, 288.05, 288.25, 288.45, 288.65, 288.85, 
    289.05, 289.25, 289.45,
  284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 285.55, 285.75, 
    285.95, 286.15, 286.35, 286.55, 286.75, 286.95, 287.15, 287.35, 287.55, 
    287.75, 287.95, 288.15, 288.35, 288.55, 288.75, 288.95, 289.15, 289.35, 
    289.55, 289.75, 289.95,
  284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 286.05, 286.25, 
    286.45, 286.65, 286.85, 287.05, 287.25, 287.45, 287.65, 287.85, 288.05, 
    288.25, 288.45, 288.65, 288.85, 289.05, 289.25, 289.45, 289.65, 289.85, 
    290.05, 290.25, 290.45,
  285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 286.55, 286.75, 
    286.95, 287.15, 287.35, 287.55, 287.75, 287.95, 288.15, 288.35, 288.55, 
    288.75, 288.95, 289.15, 289.35, 289.55, 289.75, 289.95, 290.15, 290.35, 
    290.55, 290.75, 290.95,
  285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 287.05, 287.25, 
    287.45, 287.65, 287.85, 288.05, 288.25, 288.45, 288.65, 288.85, 289.05, 
    289.25, 289.45, 289.65, 289.85, 290.05, 290.25, 290.45, 290.65, 290.85, 
    291.05, 291.25, 291.45,
  277.15, 277.35, 277.55, 277.75, 277.95, 278.15, 278.35, 278.55, 278.75, 
    278.95, 279.15, 279.35, 279.55, 279.75, 279.95, 280.15, 280.35, 280.55, 
    280.75, 280.95, 281.15, 281.35, 281.55, 281.75, 281.95, 282.15, 282.35, 
    282.55, 282.75, 282.95,
  277.65, 277.85, 278.05, 278.25, 278.45, 278.65, 278.85, 279.05, 279.25, 
    279.45, 279.65, 279.85, 280.05, 280.25, 280.45, 280.65, 280.85, 281.05, 
    281.25, 281.45, 281.65, 281.85, 282.05, 282.25, 282.45, 282.65, 282.85, 
    283.05, 283.25, 283.45,
  278.15, 278.35, 278.55, 278.75, 278.95, 279.15, 279.35, 279.55, 279.75, 
    279.95, 280.15, 280.35, 280.55, 280.75, 280.95, 281.15, 281.35, 281.55, 
    281.75, 281.95, 282.15, 282.35, 282.55, 282.75, 282.95, 283.15, 283.35, 
    283.55, 283.75, 283.95,
  278.65, 278.85, 279.05, 279.25, 279.45, 279.65, 279.85, 280.05, 280.25, 
    280.45, 280.65, 280.85, 281.05, 281.25, 281.45, 281.65, 281.85, 282.05, 
    282.25, 282.45, 282.65, 282.85, 283.05, 283.25, 283.45, 283.65, 283.85, 
    284.05, 284.25, 284.45,
  279.15, 279.35, 279.55, 279.75, 279.95, 280.15, 280.35, 280.55, 280.75, 
    280.95, 281.15, 281.35, 281.55, 281.75, 281.95, 282.15, 282.35, 282.55, 
    282.75, 282.95, 283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 
    284.55, 284.75, 284.95,
  279.65, 279.85, 280.05, 280.25, 280.45, 280.65, 280.85, 281.05, 281.25, 
    281.45, 281.65, 281.85, 282.05, 282.25, 282.45, 282.65, 282.85, 283.05, 
    283.25, 283.45, 283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 
    285.05, 285.25, 285.45,
  280.15, 280.35, 280.55, 280.75, 280.95, 281.15, 281.35, 281.55, 281.75, 
    281.95, 282.15, 282.35, 282.55, 282.75, 282.95, 283.15, 283.35, 283.55, 
    283.75, 283.95, 284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 
    285.55, 285.75, 285.95,
  280.65, 280.85, 281.05, 281.25, 281.45, 281.65, 281.85, 282.05, 282.25, 
    282.45, 282.65, 282.85, 283.05, 283.25, 283.45, 283.65, 283.85, 284.05, 
    284.25, 284.45, 284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 
    286.05, 286.25, 286.45,
  281.15, 281.35, 281.55, 281.75, 281.95, 282.15, 282.35, 282.55, 282.75, 
    282.95, 283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 284.55, 
    284.75, 284.95, 285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 
    286.55, 286.75, 286.95,
  281.65, 281.85, 282.05, 282.25, 282.45, 282.65, 282.85, 283.05, 283.25, 
    283.45, 283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 285.05, 
    285.25, 285.45, 285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 
    287.05, 287.25, 287.45,
  282.15, 282.35, 282.55, 282.75, 282.95, 283.15, 283.35, 283.55, 283.75, 
    283.95, 284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 285.55, 
    285.75, 285.95, 286.15, 286.35, 286.55, 286.75, 286.95, 287.15, 287.35, 
    287.55, 287.75, 287.95,
  282.65, 282.85, 283.05, 283.25, 283.45, 283.65, 283.85, 284.05, 284.25, 
    284.45, 284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 286.05, 
    286.25, 286.45, 286.65, 286.85, 287.05, 287.25, 287.45, 287.65, 287.85, 
    288.05, 288.25, 288.45,
  283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 284.55, 284.75, 
    284.95, 285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 286.55, 
    286.75, 286.95, 287.15, 287.35, 287.55, 287.75, 287.95, 288.15, 288.35, 
    288.55, 288.75, 288.95,
  283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 285.05, 285.25, 
    285.45, 285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 287.05, 
    287.25, 287.45, 287.65, 287.85, 288.05, 288.25, 288.45, 288.65, 288.85, 
    289.05, 289.25, 289.45,
  284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 285.55, 285.75, 
    285.95, 286.15, 286.35, 286.55, 286.75, 286.95, 287.15, 287.35, 287.55, 
    287.75, 287.95, 288.15, 288.35, 288.55, 288.75, 288.95, 289.15, 289.35, 
    289.55, 289.75, 289.95,
  284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 286.05, 286.25, 
    286.45, 286.65, 286.85, 287.05, 287.25, 287.45, 287.65, 287.85, 288.05, 
    288.25, 288.45, 288.65, 288.85, 289.05, 289.25, 289.45, 289.65, 289.85, 
    290.05, 290.25, 290.45,
  285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 286.55, 286.75, 
    286.95, 287.15, 287.35, 287.55, 287.75, 287.95, 288.15, 288.35, 288.55, 
    288.75, 288.95, 289.15, 289.35, 289.55, 289.75, 289.95, 290.15, 290.35, 
    290.55, 290.75, 290.95,
  285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 287.05, 287.25, 
    287.45, 287.65, 287.85, 288.05, 288.25, 288.45, 288.65, 288.85, 289.05, 
    289.25, 289.45, 289.65, 289.85, 290.05, 290.25, 290.45, 290.65, 290.85, 
    291.05, 291.25, 291.45,
  286.15, 286.35, 286.55, 286.75, 286.95, 287.15, 287.35, 287.55, 287.75, 
    287.95, 288.15, 288.35, 288.55, 288.75, 288.95, 289.15, 289.35, 289.55, 
    289.75, 289.95, 290.15, 290.35, 290.55, 290.75, 290.95, 291.15, 291.35, 
    291.55, 291.75, 291.95,
  286.65, 286.85, 287.05, 287.25, 287.45, 287.65, 287.85, 288.05, 288.25, 
    288.45, 288.65, 288.85, 289.05, 289.25, 289.45, 289.65, 289.85, 290.05, 
    290.25, 290.45, 290.65, 290.85, 291.05, 291.25, 291.45, 291.65, 291.85, 
    292.05, 292.25, 292.45,
  278.15, 278.35, 278.55, 278.75, 278.95, 279.15, 279.35, 279.55, 279.75, 
    279.95, 280.15, 280.35, 280.55, 280.75, 280.95, 281.15, 281.35, 281.55, 
    281.75, 281.95, 282.15, 282.35, 282.55, 282.75, 282.95, 283.15, 283.35, 
    283.55, 283.75, 283.95,
  278.65, 278.85, 279.05, 279.25, 279.45, 279.65, 279.85, 280.05, 280.25, 
    280.45, 280.65, 280.85, 281.05, 281.25, 281.45, 281.65, 281.85, 282.05, 
    282.25, 282.45, 282.65, 282.85, 283.05, 283.25, 283.45, 283.65, 283.85, 
    284.05, 284.25, 284.45,
  279.15, 279.35, 279.55, 279.75, 279.95, 280.15, 280.35, 280.55, 280.75, 
    280.95, 281.15, 281.35, 281.55, 281.75, 281.95, 282.15, 282.35, 282.55, 
    282.75, 282.95, 283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 
    284.55, 284.75, 284.95,
  279.65, 279.85, 280.05, 280.25, 280.45, 280.65, 280.85, 281.05, 281.25, 
    281.45, 281.65, 281.85, 282.05, 282.25, 282.45, 282.65, 282.85, 283.05, 
    283.25, 283.45, 283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 
    285.05, 285.25, 285.45,
  280.15, 280.35, 280.55, 280.75, 280.95, 281.15, 281.35, 281.55, 281.75, 
    281.95, 282.15, 282.35, 282.55, 282.75, 282.95, 283.15, 283.35, 283.55, 
    283.75, 283.95, 284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 
    285.55, 285.75, 285.95,
  280.65, 280.85, 281.05, 281.25, 281.45, 281.65, 281.85, 282.05, 282.25, 
    282.45, 282.65, 282.85, 283.05, 283.25, 283.45, 283.65, 283.85, 284.05, 
    284.25, 284.45, 284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 
    286.05, 286.25, 286.45,
  281.15, 281.35, 281.55, 281.75, 281.95, 282.15, 282.35, 282.55, 282.75, 
    282.95, 283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 284.55, 
    284.75, 284.95, 285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 
    286.55, 286.75, 286.95,
  281.65, 281.85, 282.05, 282.25, 282.45, 282.65, 282.85, 283.05, 283.25, 
    283.45, 283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 285.05, 
    285.25, 285.45, 285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 
    287.05, 287.25, 287.45,
  282.15, 282.35, 282.55, 282.75, 282.95, 283.15, 283.35, 283.55, 283.75, 
    283.95, 284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 285.55, 
    285.75, 285.95, 286.15, 286.35, 286.55, 286.75, 286.95, 287.15, 287.35, 
    287.55, 287.75, 287.95,
  282.65, 282.85, 283.05, 283.25, 283.45, 283.65, 283.85, 284.05, 284.25, 
    284.45, 284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 286.05, 
    286.25, 286.45, 286.65, 286.85, 287.05, 287.25, 287.45, 287.65, 287.85, 
    288.05, 288.25, 288.45,
  283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 284.55, 284.75, 
    284.95, 285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 286.55, 
    286.75, 286.95, 287.15, 287.35, 287.55, 287.75, 287.95, 288.15, 288.35, 
    288.55, 288.75, 288.95,
  283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 285.05, 285.25, 
    285.45, 285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 287.05, 
    287.25, 287.45, 287.65, 287.85, 288.05, 288.25, 288.45, 288.65, 288.85, 
    289.05, 289.25, 289.45,
  284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 285.55, 285.75, 
    285.95, 286.15, 286.35, 286.55, 286.75, 286.95, 287.15, 287.35, 287.55, 
    287.75, 287.95, 288.15, 288.35, 288.55, 288.75, 288.95, 289.15, 289.35, 
    289.55, 289.75, 289.95,
  284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 286.05, 286.25, 
    286.45, 286.65, 286.85, 287.05, 287.25, 287.45, 287.65, 287.85, 288.05, 
    288.25, 288.45, 288.65, 288.85, 289.05, 289.25, 289.45, 289.65, 289.85, 
    290.05, 290.25, 290.45,
  285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 286.55, 286.75, 
    286.95, 287.15, 287.35, 287.55, 287.75, 287.95, 288.15, 288.35, 288.55, 
    288.75, 288.95, 289.15, 289.35, 289.55, 289.75, 289.95, 290.15, 290.35, 
    290.55, 290.75, 290.95,
  285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 287.05, 287.25, 
    287.45, 287.65, 287.85, 288.05, 288.25, 288.45, 288.65, 288.85, 289.05, 
    289.25, 289.45, 289.65, 289.85, 290.05, 290.25, 290.45, 290.65, 290.85, 
    291.05, 291.25, 291.45,
  286.15, 286.35, 286.55, 286.75, 286.95, 287.15, 287.35, 287.55, 287.75, 
    287.95, 288.15, 288.35, 288.55, 288.75, 288.95, 289.15, 289.35, 289.55, 
    289.75, 289.95, 290.15, 290.35, 290.55, 290.75, 290.95, 291.15, 291.35, 
    291.55, 291.75, 291.95,
  286.65, 286.85, 287.05, 287.25, 287.45, 287.65, 287.85, 288.05, 288.25, 
    288.45, 288.65, 288.85, 289.05, 289.25, 289.45, 289.65, 289.85, 290.05, 
    290.25, 290.45, 290.65, 290.85, 291.05, 291.25, 291.45, 291.65, 291.85, 
    292.05, 292.25, 292.45,
  287.15, 287.35, 287.55, 287.75, 287.95, 288.15, 288.35, 288.55, 288.75, 
    288.95, 289.15, 289.35, 289.55, 289.75, 289.95, 290.15, 290.35, 290.55, 
    290.75, 290.95, 291.15, 291.35, 291.55, 291.75, 291.95, 292.15, 292.35, 
    292.55, 292.75, 292.95,
  287.65, 287.85, 288.05, 288.25, 288.45, 288.65, 288.85, 289.05, 289.25, 
    289.45, 289.65, 289.85, 290.05, 290.25, 290.45, 290.65, 290.85, 291.05, 
    291.25, 291.45, 291.65, 291.85, 292.05, 292.25, 292.45, 292.65, 292.85, 
    293.05, 293.25, 293.45,
  279.15, 279.35, 279.55, 279.75, 279.95, 280.15, 280.35, 280.55, 280.75, 
    280.95, 281.15, 281.35, 281.55, 281.75, 281.95, 282.15, 282.35, 282.55, 
    282.75, 282.95, 283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 
    284.55, 284.75, 284.95,
  279.65, 279.85, 280.05, 280.25, 280.45, 280.65, 280.85, 281.05, 281.25, 
    281.45, 281.65, 281.85, 282.05, 282.25, 282.45, 282.65, 282.85, 283.05, 
    283.25, 283.45, 283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 
    285.05, 285.25, 285.45,
  280.15, 280.35, 280.55, 280.75, 280.95, 281.15, 281.35, 281.55, 281.75, 
    281.95, 282.15, 282.35, 282.55, 282.75, 282.95, 283.15, 283.35, 283.55, 
    283.75, 283.95, 284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 
    285.55, 285.75, 285.95,
  280.65, 280.85, 281.05, 281.25, 281.45, 281.65, 281.85, 282.05, 282.25, 
    282.45, 282.65, 282.85, 283.05, 283.25, 283.45, 283.65, 283.85, 284.05, 
    284.25, 284.45, 284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 
    286.05, 286.25, 286.45,
  281.15, 281.35, 281.55, 281.75, 281.95, 282.15, 282.35, 282.55, 282.75, 
    282.95, 283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 284.55, 
    284.75, 284.95, 285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 
    286.55, 286.75, 286.95,
  281.65, 281.85, 282.05, 282.25, 282.45, 282.65, 282.85, 283.05, 283.25, 
    283.45, 283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 285.05, 
    285.25, 285.45, 285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 
    287.05, 287.25, 287.45,
  282.15, 282.35, 282.55, 282.75, 282.95, 283.15, 283.35, 283.55, 283.75, 
    283.95, 284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 285.55, 
    285.75, 285.95, 286.15, 286.35, 286.55, 286.75, 286.95, 287.15, 287.35, 
    287.55, 287.75, 287.95,
  282.65, 282.85, 283.05, 283.25, 283.45, 283.65, 283.85, 284.05, 284.25, 
    284.45, 284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 286.05, 
    286.25, 286.45, 286.65, 286.85, 287.05, 287.25, 287.45, 287.65, 287.85, 
    288.05, 288.25, 288.45,
  283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 284.55, 284.75, 
    284.95, 285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 286.55, 
    286.75, 286.95, 287.15, 287.35, 287.55, 287.75, 287.95, 288.15, 288.35, 
    288.55, 288.75, 288.95,
  283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 285.05, 285.25, 
    285.45, 285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 287.05, 
    287.25, 287.45, 287.65, 287.85, 288.05, 288.25, 288.45, 288.65, 288.85, 
    289.05, 289.25, 289.45,
  284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 285.55, 285.75, 
    285.95, 286.15, 286.35, 286.55, 286.75, 286.95, 287.15, 287.35, 287.55, 
    287.75, 287.95, 288.15, 288.35, 288.55, 288.75, 288.95, 289.15, 289.35, 
    289.55, 289.75, 289.95,
  284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 286.05, 286.25, 
    286.45, 286.65, 286.85, 287.05, 287.25, 287.45, 287.65, 287.85, 288.05, 
    288.25, 288.45, 288.65, 288.85, 289.05, 289.25, 289.45, 289.65, 289.85, 
    290.05, 290.25, 290.45,
  285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 286.55, 286.75, 
    286.95, 287.15, 287.35, 287.55, 287.75, 287.95, 288.15, 288.35, 288.55, 
    288.75, 288.95, 289.15, 289.35, 289.55, 289.75, 289.95, 290.15, 290.35, 
    290.55, 290.75, 290.95,
  285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 287.05, 287.25, 
    287.45, 287.65, 287.85, 288.05, 288.25, 288.45, 288.65, 288.85, 289.05, 
    289.25, 289.45, 289.65, 289.85, 290.05, 290.25, 290.45, 290.65, 290.85, 
    291.05, 291.25, 291.45,
  286.15, 286.35, 286.55, 286.75, 286.95, 287.15, 287.35, 287.55, 287.75, 
    287.95, 288.15, 288.35, 288.55, 288.75, 288.95, 289.15, 289.35, 289.55, 
    289.75, 289.95, 290.15, 290.35, 290.55, 290.75, 290.95, 291.15, 291.35, 
    291.55, 291.75, 291.95,
  286.65, 286.85, 287.05, 287.25, 287.45, 287.65, 287.85, 288.05, 288.25, 
    288.45, 288.65, 288.85, 289.05, 289.25, 289.45, 289.65, 289.85, 290.05, 
    290.25, 290.45, 290.65, 290.85, 291.05, 291.25, 291.45, 291.65, 291.85, 
    292.05, 292.25, 292.45,
  287.15, 287.35, 287.55, 287.75, 287.95, 288.15, 288.35, 288.55, 288.75, 
    288.95, 289.15, 289.35, 289.55, 289.75, 289.95, 290.15, 290.35, 290.55, 
    290.75, 290.95, 291.15, 291.35, 291.55, 291.75, 291.95, 292.15, 292.35, 
    292.55, 292.75, 292.95,
  287.65, 287.85, 288.05, 288.25, 288.45, 288.65, 288.85, 289.05, 289.25, 
    289.45, 289.65, 289.85, 290.05, 290.25, 290.45, 290.65, 290.85, 291.05, 
    291.25, 291.45, 291.65, 291.85, 292.05, 292.25, 292.45, 292.65, 292.85, 
    293.05, 293.25, 293.45,
  288.15, 288.35, 288.55, 288.75, 288.95, 289.15, 289.35, 289.55, 289.75, 
    289.95, 290.15, 290.35, 290.55, 290.75, 290.95, 291.15, 291.35, 291.55, 
    291.75, 291.95, 292.15, 292.35, 292.55, 292.75, 292.95, 293.15, 293.35, 
    293.55, 293.75, 293.95,
  288.65, 288.85, 289.05, 289.25, 289.45, 289.65, 289.85, 290.05, 290.25, 
    290.45, 290.65, 290.85, 291.05, 291.25, 291.45, 291.65, 291.85, 292.05, 
    292.25, 292.45, 292.65, 292.85, 293.05, 293.25, 293.45, 293.65, 293.85, 
    294.05, 294.25, 294.45,
  280.15, 280.35, 280.55, 280.75, 280.95, 281.15, 281.35, 281.55, 281.75, 
    281.95, 282.15, 282.35, 282.55, 282.75, 282.95, 283.15, 283.35, 283.55, 
    283.75, 283.95, 284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 
    285.55, 285.75, 285.95,
  280.65, 280.85, 281.05, 281.25, 281.45, 281.65, 281.85, 282.05, 282.25, 
    282.45, 282.65, 282.85, 283.05, 283.25, 283.45, 283.65, 283.85, 284.05, 
    284.25, 284.45, 284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 
    286.05, 286.25, 286.45,
  281.15, 281.35, 281.55, 281.75, 281.95, 282.15, 282.35, 282.55, 282.75, 
    282.95, 283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 284.55, 
    284.75, 284.95, 285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 
    286.55, 286.75, 286.95,
  281.65, 281.85, 282.05, 282.25, 282.45, 282.65, 282.85, 283.05, 283.25, 
    283.45, 283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 285.05, 
    285.25, 285.45, 285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 
    287.05, 287.25, 287.45,
  282.15, 282.35, 282.55, 282.75, 282.95, 283.15, 283.35, 283.55, 283.75, 
    283.95, 284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 285.55, 
    285.75, 285.95, 286.15, 286.35, 286.55, 286.75, 286.95, 287.15, 287.35, 
    287.55, 287.75, 287.95,
  282.65, 282.85, 283.05, 283.25, 283.45, 283.65, 283.85, 284.05, 284.25, 
    284.45, 284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 286.05, 
    286.25, 286.45, 286.65, 286.85, 287.05, 287.25, 287.45, 287.65, 287.85, 
    288.05, 288.25, 288.45,
  283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 284.55, 284.75, 
    284.95, 285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 286.55, 
    286.75, 286.95, 287.15, 287.35, 287.55, 287.75, 287.95, 288.15, 288.35, 
    288.55, 288.75, 288.95,
  283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 285.05, 285.25, 
    285.45, 285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 287.05, 
    287.25, 287.45, 287.65, 287.85, 288.05, 288.25, 288.45, 288.65, 288.85, 
    289.05, 289.25, 289.45,
  284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 285.55, 285.75, 
    285.95, 286.15, 286.35, 286.55, 286.75, 286.95, 287.15, 287.35, 287.55, 
    287.75, 287.95, 288.15, 288.35, 288.55, 288.75, 288.95, 289.15, 289.35, 
    289.55, 289.75, 289.95,
  284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 286.05, 286.25, 
    286.45, 286.65, 286.85, 287.05, 287.25, 287.45, 287.65, 287.85, 288.05, 
    288.25, 288.45, 288.65, 288.85, 289.05, 289.25, 289.45, 289.65, 289.85, 
    290.05, 290.25, 290.45,
  285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 286.55, 286.75, 
    286.95, 287.15, 287.35, 287.55, 287.75, 287.95, 288.15, 288.35, 288.55, 
    288.75, 288.95, 289.15, 289.35, 289.55, 289.75, 289.95, 290.15, 290.35, 
    290.55, 290.75, 290.95,
  285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 287.05, 287.25, 
    287.45, 287.65, 287.85, 288.05, 288.25, 288.45, 288.65, 288.85, 289.05, 
    289.25, 289.45, 289.65, 289.85, 290.05, 290.25, 290.45, 290.65, 290.85, 
    291.05, 291.25, 291.45,
  286.15, 286.35, 286.55, 286.75, 286.95, 287.15, 287.35, 287.55, 287.75, 
    287.95, 288.15, 288.35, 288.55, 288.75, 288.95, 289.15, 289.35, 289.55, 
    289.75, 289.95, 290.15, 290.35, 290.55, 290.75, 290.95, 291.15, 291.35, 
    291.55, 291.75, 291.95,
  286.65, 286.85, 287.05, 287.25, 287.45, 287.65, 287.85, 288.05, 288.25, 
    288.45, 288.65, 288.85, 289.05, 289.25, 289.45, 289.65, 289.85, 290.05, 
    290.25, 290.45, 290.65, 290.85, 291.05, 291.25, 291.45, 291.65, 291.85, 
    292.05, 292.25, 292.45,
  287.15, 287.35, 287.55, 287.75, 287.95, 288.15, 288.35, 288.55, 288.75, 
    288.95, 289.15, 289.35, 289.55, 289.75, 289.95, 290.15, 290.35, 290.55, 
    290.75, 290.95, 291.15, 291.35, 291.55, 291.75, 291.95, 292.15, 292.35, 
    292.55, 292.75, 292.95,
  287.65, 287.85, 288.05, 288.25, 288.45, 288.65, 288.85, 289.05, 289.25, 
    289.45, 289.65, 289.85, 290.05, 290.25, 290.45, 290.65, 290.85, 291.05, 
    291.25, 291.45, 291.65, 291.85, 292.05, 292.25, 292.45, 292.65, 292.85, 
    293.05, 293.25, 293.45,
  288.15, 288.35, 288.55, 288.75, 288.95, 289.15, 289.35, 289.55, 289.75, 
    289.95, 290.15, 290.35, 290.55, 290.75, 290.95, 291.15, 291.35, 291.55, 
    291.75, 291.95, 292.15, 292.35, 292.55, 292.75, 292.95, 293.15, 293.35, 
    293.55, 293.75, 293.95,
  288.65, 288.85, 289.05, 289.25, 289.45, 289.65, 289.85, 290.05, 290.25, 
    290.45, 290.65, 290.85, 291.05, 291.25, 291.45, 291.65, 291.85, 292.05, 
    292.25, 292.45, 292.65, 292.85, 293.05, 293.25, 293.45, 293.65, 293.85, 
    294.05, 294.25, 294.45,
  289.15, 289.35, 289.55, 289.75, 289.95, 290.15, 290.35, 290.55, 290.75, 
    290.95, 291.15, 291.35, 291.55, 291.75, 291.95, 292.15, 292.35, 292.55, 
    292.75, 292.95, 293.15, 293.35, 293.55, 293.75, 293.95, 294.15, 294.35, 
    294.55, 294.75, 294.95,
  289.65, 289.85, 290.05, 290.25, 290.45, 290.65, 290.85, 291.05, 291.25, 
    291.45, 291.65, 291.85, 292.05, 292.25, 292.45, 292.65, 292.85, 293.05, 
    293.25, 293.45, 293.65, 293.85, 294.05, 294.25, 294.45, 294.65, 294.85, 
    295.05, 295.25, 295.45,
  281.15, 281.35, 281.55, 281.75, 281.95, 282.15, 282.35, 282.55, 282.75, 
    282.95, 283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 284.55, 
    284.75, 284.95, 285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 
    286.55, 286.75, 286.95,
  281.65, 281.85, 282.05, 282.25, 282.45, 282.65, 282.85, 283.05, 283.25, 
    283.45, 283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 285.05, 
    285.25, 285.45, 285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 
    287.05, 287.25, 287.45,
  282.15, 282.35, 282.55, 282.75, 282.95, 283.15, 283.35, 283.55, 283.75, 
    283.95, 284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 285.55, 
    285.75, 285.95, 286.15, 286.35, 286.55, 286.75, 286.95, 287.15, 287.35, 
    287.55, 287.75, 287.95,
  282.65, 282.85, 283.05, 283.25, 283.45, 283.65, 283.85, 284.05, 284.25, 
    284.45, 284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 286.05, 
    286.25, 286.45, 286.65, 286.85, 287.05, 287.25, 287.45, 287.65, 287.85, 
    288.05, 288.25, 288.45,
  283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 284.55, 284.75, 
    284.95, 285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 286.55, 
    286.75, 286.95, 287.15, 287.35, 287.55, 287.75, 287.95, 288.15, 288.35, 
    288.55, 288.75, 288.95,
  283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 285.05, 285.25, 
    285.45, 285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 287.05, 
    287.25, 287.45, 287.65, 287.85, 288.05, 288.25, 288.45, 288.65, 288.85, 
    289.05, 289.25, 289.45,
  284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 285.55, 285.75, 
    285.95, 286.15, 286.35, 286.55, 286.75, 286.95, 287.15, 287.35, 287.55, 
    287.75, 287.95, 288.15, 288.35, 288.55, 288.75, 288.95, 289.15, 289.35, 
    289.55, 289.75, 289.95,
  284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 286.05, 286.25, 
    286.45, 286.65, 286.85, 287.05, 287.25, 287.45, 287.65, 287.85, 288.05, 
    288.25, 288.45, 288.65, 288.85, 289.05, 289.25, 289.45, 289.65, 289.85, 
    290.05, 290.25, 290.45,
  285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 286.55, 286.75, 
    286.95, 287.15, 287.35, 287.55, 287.75, 287.95, 288.15, 288.35, 288.55, 
    288.75, 288.95, 289.15, 289.35, 289.55, 289.75, 289.95, 290.15, 290.35, 
    290.55, 290.75, 290.95,
  285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 287.05, 287.25, 
    287.45, 287.65, 287.85, 288.05, 288.25, 288.45, 288.65, 288.85, 289.05, 
    289.25, 289.45, 289.65, 289.85, 290.05, 290.25, 290.45, 290.65, 290.85, 
    291.05, 291.25, 291.45,
  286.15, 286.35, 286.55, 286.75, 286.95, 287.15, 287.35, 287.55, 287.75, 
    287.95, 288.15, 288.35, 288.55, 288.75, 288.95, 289.15, 289.35, 289.55, 
    289.75, 289.95, 290.15, 290.35, 290.55, 290.75, 290.95, 291.15, 291.35, 
    291.55, 291.75, 291.95,
  286.65, 286.85, 287.05, 287.25, 287.45, 287.65, 287.85, 288.05, 288.25, 
    288.45, 288.65, 288.85, 289.05, 289.25, 289.45, 289.65, 289.85, 290.05, 
    290.25, 290.45, 290.65, 290.85, 291.05, 291.25, 291.45, 291.65, 291.85, 
    292.05, 292.25, 292.45,
  287.15, 287.35, 287.55, 287.75, 287.95, 288.15, 288.35, 288.55, 288.75, 
    288.95, 289.15, 289.35, 289.55, 289.75, 289.95, 290.15, 290.35, 290.55, 
    290.75, 290.95, 291.15, 291.35, 291.55, 291.75, 291.95, 292.15, 292.35, 
    292.55, 292.75, 292.95,
  287.65, 287.85, 288.05, 288.25, 288.45, 288.65, 288.85, 289.05, 289.25, 
    289.45, 289.65, 289.85, 290.05, 290.25, 290.45, 290.65, 290.85, 291.05, 
    291.25, 291.45, 291.65, 291.85, 292.05, 292.25, 292.45, 292.65, 292.85, 
    293.05, 293.25, 293.45,
  288.15, 288.35, 288.55, 288.75, 288.95, 289.15, 289.35, 289.55, 289.75, 
    289.95, 290.15, 290.35, 290.55, 290.75, 290.95, 291.15, 291.35, 291.55, 
    291.75, 291.95, 292.15, 292.35, 292.55, 292.75, 292.95, 293.15, 293.35, 
    293.55, 293.75, 293.95,
  288.65, 288.85, 289.05, 289.25, 289.45, 289.65, 289.85, 290.05, 290.25, 
    290.45, 290.65, 290.85, 291.05, 291.25, 291.45, 291.65, 291.85, 292.05, 
    292.25, 292.45, 292.65, 292.85, 293.05, 293.25, 293.45, 293.65, 293.85, 
    294.05, 294.25, 294.45,
  289.15, 289.35, 289.55, 289.75, 289.95, 290.15, 290.35, 290.55, 290.75, 
    290.95, 291.15, 291.35, 291.55, 291.75, 291.95, 292.15, 292.35, 292.55, 
    292.75, 292.95, 293.15, 293.35, 293.55, 293.75, 293.95, 294.15, 294.35, 
    294.55, 294.75, 294.95,
  289.65, 289.85, 290.05, 290.25, 290.45, 290.65, 290.85, 291.05, 291.25, 
    291.45, 291.65, 291.85, 292.05, 292.25, 292.45, 292.65, 292.85, 293.05, 
    293.25, 293.45, 293.65, 293.85, 294.05, 294.25, 294.45, 294.65, 294.85, 
    295.05, 295.25, 295.45,
  290.15, 290.35, 290.55, 290.75, 290.95, 291.15, 291.35, 291.55, 291.75, 
    291.95, 292.15, 292.35, 292.55, 292.75, 292.95, 293.15, 293.35, 293.55, 
    293.75, 293.95, 294.15, 294.35, 294.55, 294.75, 294.95, 295.15, 295.35, 
    295.55, 295.75, 295.95,
  290.65, 290.85, 291.05, 291.25, 291.45, 291.65, 291.85, 292.05, 292.25, 
    292.45, 292.65, 292.85, 293.05, 293.25, 293.45, 293.65, 293.85, 294.05, 
    294.25, 294.45, 294.65, 294.85, 295.05, 295.25, 295.45, 295.65, 295.85, 
    296.05, 296.25, 296.45,
  282.15, 282.35, 282.55, 282.75, 282.95, 283.15, 283.35, 283.55, 283.75, 
    283.95, 284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 285.55, 
    285.75, 285.95, 286.15, 286.35, 286.55, 286.75, 286.95, 287.15, 287.35, 
    287.55, 287.75, 287.95,
  282.65, 282.85, 283.05, 283.25, 283.45, 283.65, 283.85, 284.05, 284.25, 
    284.45, 284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 286.05, 
    286.25, 286.45, 286.65, 286.85, 287.05, 287.25, 287.45, 287.65, 287.85, 
    288.05, 288.25, 288.45,
  283.15, 283.35, 283.55, 283.75, 283.95, 284.15, 284.35, 284.55, 284.75, 
    284.95, 285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 286.55, 
    286.75, 286.95, 287.15, 287.35, 287.55, 287.75, 287.95, 288.15, 288.35, 
    288.55, 288.75, 288.95,
  283.65, 283.85, 284.05, 284.25, 284.45, 284.65, 284.85, 285.05, 285.25, 
    285.45, 285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 287.05, 
    287.25, 287.45, 287.65, 287.85, 288.05, 288.25, 288.45, 288.65, 288.85, 
    289.05, 289.25, 289.45,
  284.15, 284.35, 284.55, 284.75, 284.95, 285.15, 285.35, 285.55, 285.75, 
    285.95, 286.15, 286.35, 286.55, 286.75, 286.95, 287.15, 287.35, 287.55, 
    287.75, 287.95, 288.15, 288.35, 288.55, 288.75, 288.95, 289.15, 289.35, 
    289.55, 289.75, 289.95,
  284.65, 284.85, 285.05, 285.25, 285.45, 285.65, 285.85, 286.05, 286.25, 
    286.45, 286.65, 286.85, 287.05, 287.25, 287.45, 287.65, 287.85, 288.05, 
    288.25, 288.45, 288.65, 288.85, 289.05, 289.25, 289.45, 289.65, 289.85, 
    290.05, 290.25, 290.45,
  285.15, 285.35, 285.55, 285.75, 285.95, 286.15, 286.35, 286.55, 286.75, 
    286.95, 287.15, 287.35, 287.55, 287.75, 287.95, 288.15, 288.35, 288.55, 
    288.75, 288.95, 289.15, 289.35, 289.55, 289.75, 289.95, 290.15, 290.35, 
    290.55, 290.75, 290.95,
  285.65, 285.85, 286.05, 286.25, 286.45, 286.65, 286.85, 287.05, 287.25, 
    287.45, 287.65, 287.85, 288.05, 288.25, 288.45, 288.65, 288.85, 289.05, 
    289.25, 289.45, 289.65, 289.85, 290.05, 290.25, 290.45, 290.65, 290.85, 
    291.05, 291.25, 291.45,
  286.15, 286.35, 286.55, 286.75, 286.95, 287.15, 287.35, 287.55, 287.75, 
    287.95, 288.15, 288.35, 288.55, 288.75, 288.95, 289.15, 289.35, 289.55, 
    289.75, 289.95, 290.15, 290.35, 290.55, 290.75, 290.95, 291.15, 291.35, 
    291.55, 291.75, 291.95,
  286.65, 286.85, 287.05, 287.25, 287.45, 287.65, 287.85, 288.05, 288.25, 
    288.45, 288.65, 288.85, 289.05, 289.25, 289.45, 289.65, 289.85, 290.05, 
    290.25, 290.45, 290.65, 290.85, 291.05, 291.25, 291.45, 291.65, 291.85, 
    292.05, 292.25, 292.45,
  287.15, 287.35, 287.55, 287.75, 287.95, 288.15, 288.35, 288.55, 288.75, 
    288.95, 289.15, 289.35, 289.55, 289.75, 289.95, 290.15, 290.35, 290.55, 
    290.75, 290.95, 291.15, 291.35, 291.55, 291.75, 291.95, 292.15, 292.35, 
    292.55, 292.75, 292.95,
  287.65, 287.85, 288.05, 288.25, 288.45, 288.65, 288.85, 289.05, 289.25, 
    289.45, 289.65, 289.85, 290.05, 290.25, 290.45, 290.65, 290.85, 291.05, 
    291.25, 291.45, 291.65, 291.85, 292.05, 292.25, 292.45, 292.65, 292.85, 
    293.05, 293.25, 293.45,
  288.15, 288.35, 288.55, 288.75, 288.95, 289.15, 289.35, 289.55, 289.75, 
    289.95, 290.15, 290.35, 290.55, 290.75, 290.95, 291.15, 291.35, 291.55, 
    291.75, 291.95, 292.15, 292.35, 292.55, 292.75, 292.95, 293.15, 293.35, 
    293.55, 293.75, 293.95,
  288.65, 288.85, 289.05, 289.25, 289.45, 289.65, 289.85, 290.05, 290.25, 
    290.45, 290.65, 290.85, 291.05, 291.25, 291.45, 291.65, 291.85, 292.05, 
    292.25, 292.45, 292.65, 292.85, 293.05, 293.25, 293.45, 293.65, 293.85, 
    294.05, 294.25, 294.45,
  289.15, 289.35, 289.55, 289.75, 289.95, 290.15, 290.35, 290.55, 290.75, 
    290.95, 291.15, 291.35, 291.55, 291.75, 291.95, 292.15, 292.35, 292.55, 
    292.75, 292.95, 293.15, 293.35, 293.55, 293.75, 293.95, 294.15, 294.35, 
    294.55, 294.75, 294.95,
  289.65, 289.85, 290.05, 290.25, 290.45, 290.65, 290.85, 291.05, 291.25, 
    291.45, 291.65, 291.85, 292.05, 292.25, 292.45, 292.65, 292.85, 293.05, 
    293.25, 293.45, 293.65, 293.85, 294.05, 294.25, 294.45, 294.65, 294.85, 
    295.05, 295.25, 295.45,
  290.15, 290.35, 290.55, 290.75, 290.95, 291.15, 291.35, 291.55, 291.75, 
    291.95, 292.15, 292.35, 292.55, 292.75, 292.95, 293.15, 293.35, 293.55, 
    293.75, 293.95, 294.15, 294.35, 294.55, 294.75, 294.95, 295.15, 295.35, 
    295.55, 295.75, 295.95,
  290.65, 290.85, 291.05, 291.25, 291.45, 291.65, 291.85, 292.05, 292.25, 
    292.45, 292.65, 292.85, 293.05, 293.25, 293.45, 293.65, 293.85, 294.05, 
    294.25, 294.45, 294.65, 294.85, 295.05, 295.25, 295.45, 295.65, 295.85, 
    296.05, 296.25, 296.45,
  291.15, 291.35, 291.55, 291.75, 291.95, 292.15, 292.35, 292.55, 292.75, 
    292.95, 293.15, 293.35, 293.55, 293.75, 293.95, 294.15, 294.35, 294.55, 
    294.75, 294.95, 295.15, 295.35, 295.55, 295.75, 295.95, 296.15, 296.35, 
    296.55, 296.75, 296.95,
  291.65, 291.85, 292.05, 292.25, 292.45, 292.65, 292.85, 293.05, 293.25, 
    293.45, 293.65, 293.85, 294.05, 294.25, 294.45, 294.65, 294.85, 295.05, 
    295.25, 295.45, 295.65, 295.85, 296.05, 296.25, 296.45, 296.65, 296.85, 
    297.05, 297.25, 297.45 ;

 pressure =
  1013.25, 1013.27, 1013.29, 1013.31, 1013.33, 1013.35, 1013.37, 1013.39, 
    1013.41, 1013.43, 1013.45, 1013.47, 1013.49, 1013.51, 1013.53, 1013.55, 
    1013.57, 1013.59, 1013.61, 1013.63, 1013.65, 1013.67, 1013.69, 1013.71, 
    1013.73, 1013.75, 1013.77, 1013.79, 1013.81, 1013.83,
  1013.3, 1013.32, 1013.34, 1013.36, 1013.38, 1013.4, 1013.42, 1013.44, 
    1013.46, 1013.48, 1013.5, 1013.52, 1013.54, 1013.56, 1013.58, 1013.6, 
    1013.62, 1013.64, 1013.66, 1013.68, 1013.7, 1013.72, 1013.74, 1013.76, 
    1013.78, 1013.8, 1013.82, 1013.84, 1013.86, 1013.88,
  1013.35, 1013.37, 1013.39, 1013.41, 1013.43, 1013.45, 1013.47, 1013.49, 
    1013.51, 1013.53, 1013.55, 1013.57, 1013.59, 1013.61, 1013.63, 1013.65, 
    1013.67, 1013.69, 1013.71, 1013.73, 1013.75, 1013.77, 1013.79, 1013.81, 
    1013.83, 1013.85, 1013.87, 1013.89, 1013.91, 1013.93,
  1013.4, 1013.42, 1013.44, 1013.46, 1013.48, 1013.5, 1013.52, 1013.54, 
    1013.56, 1013.58, 1013.6, 1013.62, 1013.64, 1013.66, 1013.68, 1013.7, 
    1013.72, 1013.74, 1013.76, 1013.78, 1013.8, 1013.82, 1013.84, 1013.86, 
    1013.88, 1013.9, 1013.92, 1013.94, 1013.96, 1013.98,
  1013.45, 1013.47, 1013.49, 1013.51, 1013.53, 1013.55, 1013.57, 1013.59, 
    1013.61, 1013.63, 1013.65, 1013.67, 1013.69, 1013.71, 1013.73, 1013.75, 
    1013.77, 1013.79, 1013.81, 1013.83, 1013.85, 1013.87, 1013.89, 1013.91, 
    1013.93, 1013.95, 1013.97, 1013.99, 1014.01, 1014.03,
  1013.5, 1013.52, 1013.54, 1013.56, 1013.58, 1013.6, 1013.62, 1013.64, 
    1013.66, 1013.68, 1013.7, 1013.72, 1013.74, 1013.76, 1013.78, 1013.8, 
    1013.82, 1013.84, 1013.86, 1013.88, 1013.9, 1013.92, 1013.94, 1013.96, 
    1013.98, 1014, 1014.02, 1014.04, 1014.06, 1014.08,
  1013.55, 1013.57, 1013.59, 1013.61, 1013.63, 1013.65, 1013.67, 1013.69, 
    1013.71, 1013.73, 1013.75, 1013.77, 1013.79, 1013.81, 1013.83, 1013.85, 
    1013.87, 1013.89, 1013.91, 1013.93, 1013.95, 1013.97, 1013.99, 1014.01, 
    1014.03, 1014.05, 1014.07, 1014.09, 1014.11, 1014.13,
  1013.6, 1013.62, 1013.64, 1013.66, 1013.68, 1013.7, 1013.72, 1013.74, 
    1013.76, 1013.78, 1013.8, 1013.82, 1013.84, 1013.86, 1013.88, 1013.9, 
    1013.92, 1013.94, 1013.96, 1013.98, 1014, 1014.02, 1014.04, 1014.06, 
    1014.08, 1014.1, 1014.12, 1014.14, 1014.16, 1014.18,
  1013.65, 1013.67, 1013.69, 1013.71, 1013.73, 1013.75, 1013.77, 1013.79, 
    1013.81, 1013.83, 1013.85, 1013.87, 1013.89, 1013.91, 1013.93, 1013.95, 
    1013.97, 1013.99, 1014.01, 1014.03, 1014.05, 1014.07, 1014.09, 1014.11, 
    1014.13, 1014.15, 1014.17, 1014.19, 1014.21, 1014.23,
  1013.7, 1013.72, 1013.74, 1013.76, 1013.78, 1013.8, 1013.82, 1013.84, 
    1013.86, 1013.88, 1013.9, 1013.92, 1013.94, 1013.96, 1013.98, 1014, 
    1014.02, 1014.04, 1014.06, 1014.08, 1014.1, 1014.12, 1014.14, 1014.16, 
    1014.18, 1014.2, 1014.22, 1014.24, 1014.26, 1014.28,
  1013.75, 1013.77, 1013.79, 1013.81, 1013.83, 1013.85, 1013.87, 1013.89, 
    1013.91, 1013.93, 1013.95, 1013.97, 1013.99, 1014.01, 1014.03, 1014.05, 
    1014.07, 1014.09, 1014.11, 1014.13, 1014.15, 1014.17, 1014.19, 1014.21, 
    1014.23, 1014.25, 1014.27, 1014.29, 1014.31, 1014.33,
  1013.8, 1013.82, 1013.84, 1013.86, 1013.88, 1013.9, 1013.92, 1013.94, 
    1013.96, 1013.98, 1014, 1014.02, 1014.04, 1014.06, 1014.08, 1014.1, 
    1014.12, 1014.14, 1014.16, 1014.18, 1014.2, 1014.22, 1014.24, 1014.26, 
    1014.28, 1014.3, 1014.32, 1014.34, 1014.36, 1014.38,
  1013.85, 1013.87, 1013.89, 1013.91, 1013.93, 1013.95, 1013.97, 1013.99, 
    1014.01, 1014.03, 1014.05, 1014.07, 1014.09, 1014.11, 1014.13, 1014.15, 
    1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 1014.31, 
    1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 1014.43,
  1013.9, 1013.92, 1013.94, 1013.96, 1013.98, 1014, 1014.02, 1014.04, 
    1014.06, 1014.08, 1014.1, 1014.12, 1014.14, 1014.16, 1014.18, 1014.2, 
    1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 1014.36, 
    1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 1014.48,
  1013.95, 1013.97, 1013.99, 1014.01, 1014.03, 1014.05, 1014.07, 1014.09, 
    1014.11, 1014.13, 1014.15, 1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 
    1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 
    1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 1014.53,
  1014, 1014.02, 1014.04, 1014.06, 1014.08, 1014.1, 1014.12, 1014.14, 
    1014.16, 1014.18, 1014.2, 1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 
    1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 
    1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 1014.58,
  1014.05, 1014.07, 1014.09, 1014.11, 1014.13, 1014.15, 1014.17, 1014.19, 
    1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 
    1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 
    1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 1014.63,
  1014.1, 1014.12, 1014.14, 1014.16, 1014.18, 1014.2, 1014.22, 1014.24, 
    1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 
    1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 
    1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 1014.68,
  1014.15, 1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 
    1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 
    1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 
    1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 1014.73,
  1014.2, 1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 
    1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 
    1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 
    1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 1014.78,
  1013.35, 1013.37, 1013.39, 1013.41, 1013.43, 1013.45, 1013.47, 1013.49, 
    1013.51, 1013.53, 1013.55, 1013.57, 1013.59, 1013.61, 1013.63, 1013.65, 
    1013.67, 1013.69, 1013.71, 1013.73, 1013.75, 1013.77, 1013.79, 1013.81, 
    1013.83, 1013.85, 1013.87, 1013.89, 1013.91, 1013.93,
  1013.4, 1013.42, 1013.44, 1013.46, 1013.48, 1013.5, 1013.52, 1013.54, 
    1013.56, 1013.58, 1013.6, 1013.62, 1013.64, 1013.66, 1013.68, 1013.7, 
    1013.72, 1013.74, 1013.76, 1013.78, 1013.8, 1013.82, 1013.84, 1013.86, 
    1013.88, 1013.9, 1013.92, 1013.94, 1013.96, 1013.98,
  1013.45, 1013.47, 1013.49, 1013.51, 1013.53, 1013.55, 1013.57, 1013.59, 
    1013.61, 1013.63, 1013.65, 1013.67, 1013.69, 1013.71, 1013.73, 1013.75, 
    1013.77, 1013.79, 1013.81, 1013.83, 1013.85, 1013.87, 1013.89, 1013.91, 
    1013.93, 1013.95, 1013.97, 1013.99, 1014.01, 1014.03,
  1013.5, 1013.52, 1013.54, 1013.56, 1013.58, 1013.6, 1013.62, 1013.64, 
    1013.66, 1013.68, 1013.7, 1013.72, 1013.74, 1013.76, 1013.78, 1013.8, 
    1013.82, 1013.84, 1013.86, 1013.88, 1013.9, 1013.92, 1013.94, 1013.96, 
    1013.98, 1014, 1014.02, 1014.04, 1014.06, 1014.08,
  1013.55, 1013.57, 1013.59, 1013.61, 1013.63, 1013.65, 1013.67, 1013.69, 
    1013.71, 1013.73, 1013.75, 1013.77, 1013.79, 1013.81, 1013.83, 1013.85, 
    1013.87, 1013.89, 1013.91, 1013.93, 1013.95, 1013.97, 1013.99, 1014.01, 
    1014.03, 1014.05, 1014.07, 1014.09, 1014.11, 1014.13,
  1013.6, 1013.62, 1013.64, 1013.66, 1013.68, 1013.7, 1013.72, 1013.74, 
    1013.76, 1013.78, 1013.8, 1013.82, 1013.84, 1013.86, 1013.88, 1013.9, 
    1013.92, 1013.94, 1013.96, 1013.98, 1014, 1014.02, 1014.04, 1014.06, 
    1014.08, 1014.1, 1014.12, 1014.14, 1014.16, 1014.18,
  1013.65, 1013.67, 1013.69, 1013.71, 1013.73, 1013.75, 1013.77, 1013.79, 
    1013.81, 1013.83, 1013.85, 1013.87, 1013.89, 1013.91, 1013.93, 1013.95, 
    1013.97, 1013.99, 1014.01, 1014.03, 1014.05, 1014.07, 1014.09, 1014.11, 
    1014.13, 1014.15, 1014.17, 1014.19, 1014.21, 1014.23,
  1013.7, 1013.72, 1013.74, 1013.76, 1013.78, 1013.8, 1013.82, 1013.84, 
    1013.86, 1013.88, 1013.9, 1013.92, 1013.94, 1013.96, 1013.98, 1014, 
    1014.02, 1014.04, 1014.06, 1014.08, 1014.1, 1014.12, 1014.14, 1014.16, 
    1014.18, 1014.2, 1014.22, 1014.24, 1014.26, 1014.28,
  1013.75, 1013.77, 1013.79, 1013.81, 1013.83, 1013.85, 1013.87, 1013.89, 
    1013.91, 1013.93, 1013.95, 1013.97, 1013.99, 1014.01, 1014.03, 1014.05, 
    1014.07, 1014.09, 1014.11, 1014.13, 1014.15, 1014.17, 1014.19, 1014.21, 
    1014.23, 1014.25, 1014.27, 1014.29, 1014.31, 1014.33,
  1013.8, 1013.82, 1013.84, 1013.86, 1013.88, 1013.9, 1013.92, 1013.94, 
    1013.96, 1013.98, 1014, 1014.02, 1014.04, 1014.06, 1014.08, 1014.1, 
    1014.12, 1014.14, 1014.16, 1014.18, 1014.2, 1014.22, 1014.24, 1014.26, 
    1014.28, 1014.3, 1014.32, 1014.34, 1014.36, 1014.38,
  1013.85, 1013.87, 1013.89, 1013.91, 1013.93, 1013.95, 1013.97, 1013.99, 
    1014.01, 1014.03, 1014.05, 1014.07, 1014.09, 1014.11, 1014.13, 1014.15, 
    1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 1014.31, 
    1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 1014.43,
  1013.9, 1013.92, 1013.94, 1013.96, 1013.98, 1014, 1014.02, 1014.04, 
    1014.06, 1014.08, 1014.1, 1014.12, 1014.14, 1014.16, 1014.18, 1014.2, 
    1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 1014.36, 
    1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 1014.48,
  1013.95, 1013.97, 1013.99, 1014.01, 1014.03, 1014.05, 1014.07, 1014.09, 
    1014.11, 1014.13, 1014.15, 1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 
    1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 
    1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 1014.53,
  1014, 1014.02, 1014.04, 1014.06, 1014.08, 1014.1, 1014.12, 1014.14, 
    1014.16, 1014.18, 1014.2, 1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 
    1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 
    1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 1014.58,
  1014.05, 1014.07, 1014.09, 1014.11, 1014.13, 1014.15, 1014.17, 1014.19, 
    1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 
    1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 
    1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 1014.63,
  1014.1, 1014.12, 1014.14, 1014.16, 1014.18, 1014.2, 1014.22, 1014.24, 
    1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 
    1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 
    1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 1014.68,
  1014.15, 1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 
    1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 
    1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 
    1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 1014.73,
  1014.2, 1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 
    1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 
    1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 
    1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 1014.78,
  1014.25, 1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 
    1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 
    1014.57, 1014.59, 1014.61, 1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 
    1014.73, 1014.75, 1014.77, 1014.79, 1014.81, 1014.83,
  1014.3, 1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 
    1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 
    1014.62, 1014.64, 1014.66, 1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 
    1014.78, 1014.8, 1014.82, 1014.84, 1014.86, 1014.88,
  1013.45, 1013.47, 1013.49, 1013.51, 1013.53, 1013.55, 1013.57, 1013.59, 
    1013.61, 1013.63, 1013.65, 1013.67, 1013.69, 1013.71, 1013.73, 1013.75, 
    1013.77, 1013.79, 1013.81, 1013.83, 1013.85, 1013.87, 1013.89, 1013.91, 
    1013.93, 1013.95, 1013.97, 1013.99, 1014.01, 1014.03,
  1013.5, 1013.52, 1013.54, 1013.56, 1013.58, 1013.6, 1013.62, 1013.64, 
    1013.66, 1013.68, 1013.7, 1013.72, 1013.74, 1013.76, 1013.78, 1013.8, 
    1013.82, 1013.84, 1013.86, 1013.88, 1013.9, 1013.92, 1013.94, 1013.96, 
    1013.98, 1014, 1014.02, 1014.04, 1014.06, 1014.08,
  1013.55, 1013.57, 1013.59, 1013.61, 1013.63, 1013.65, 1013.67, 1013.69, 
    1013.71, 1013.73, 1013.75, 1013.77, 1013.79, 1013.81, 1013.83, 1013.85, 
    1013.87, 1013.89, 1013.91, 1013.93, 1013.95, 1013.97, 1013.99, 1014.01, 
    1014.03, 1014.05, 1014.07, 1014.09, 1014.11, 1014.13,
  1013.6, 1013.62, 1013.64, 1013.66, 1013.68, 1013.7, 1013.72, 1013.74, 
    1013.76, 1013.78, 1013.8, 1013.82, 1013.84, 1013.86, 1013.88, 1013.9, 
    1013.92, 1013.94, 1013.96, 1013.98, 1014, 1014.02, 1014.04, 1014.06, 
    1014.08, 1014.1, 1014.12, 1014.14, 1014.16, 1014.18,
  1013.65, 1013.67, 1013.69, 1013.71, 1013.73, 1013.75, 1013.77, 1013.79, 
    1013.81, 1013.83, 1013.85, 1013.87, 1013.89, 1013.91, 1013.93, 1013.95, 
    1013.97, 1013.99, 1014.01, 1014.03, 1014.05, 1014.07, 1014.09, 1014.11, 
    1014.13, 1014.15, 1014.17, 1014.19, 1014.21, 1014.23,
  1013.7, 1013.72, 1013.74, 1013.76, 1013.78, 1013.8, 1013.82, 1013.84, 
    1013.86, 1013.88, 1013.9, 1013.92, 1013.94, 1013.96, 1013.98, 1014, 
    1014.02, 1014.04, 1014.06, 1014.08, 1014.1, 1014.12, 1014.14, 1014.16, 
    1014.18, 1014.2, 1014.22, 1014.24, 1014.26, 1014.28,
  1013.75, 1013.77, 1013.79, 1013.81, 1013.83, 1013.85, 1013.87, 1013.89, 
    1013.91, 1013.93, 1013.95, 1013.97, 1013.99, 1014.01, 1014.03, 1014.05, 
    1014.07, 1014.09, 1014.11, 1014.13, 1014.15, 1014.17, 1014.19, 1014.21, 
    1014.23, 1014.25, 1014.27, 1014.29, 1014.31, 1014.33,
  1013.8, 1013.82, 1013.84, 1013.86, 1013.88, 1013.9, 1013.92, 1013.94, 
    1013.96, 1013.98, 1014, 1014.02, 1014.04, 1014.06, 1014.08, 1014.1, 
    1014.12, 1014.14, 1014.16, 1014.18, 1014.2, 1014.22, 1014.24, 1014.26, 
    1014.28, 1014.3, 1014.32, 1014.34, 1014.36, 1014.38,
  1013.85, 1013.87, 1013.89, 1013.91, 1013.93, 1013.95, 1013.97, 1013.99, 
    1014.01, 1014.03, 1014.05, 1014.07, 1014.09, 1014.11, 1014.13, 1014.15, 
    1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 1014.31, 
    1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 1014.43,
  1013.9, 1013.92, 1013.94, 1013.96, 1013.98, 1014, 1014.02, 1014.04, 
    1014.06, 1014.08, 1014.1, 1014.12, 1014.14, 1014.16, 1014.18, 1014.2, 
    1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 1014.36, 
    1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 1014.48,
  1013.95, 1013.97, 1013.99, 1014.01, 1014.03, 1014.05, 1014.07, 1014.09, 
    1014.11, 1014.13, 1014.15, 1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 
    1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 
    1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 1014.53,
  1014, 1014.02, 1014.04, 1014.06, 1014.08, 1014.1, 1014.12, 1014.14, 
    1014.16, 1014.18, 1014.2, 1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 
    1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 
    1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 1014.58,
  1014.05, 1014.07, 1014.09, 1014.11, 1014.13, 1014.15, 1014.17, 1014.19, 
    1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 
    1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 
    1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 1014.63,
  1014.1, 1014.12, 1014.14, 1014.16, 1014.18, 1014.2, 1014.22, 1014.24, 
    1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 
    1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 
    1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 1014.68,
  1014.15, 1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 
    1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 
    1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 
    1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 1014.73,
  1014.2, 1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 
    1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 
    1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 
    1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 1014.78,
  1014.25, 1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 
    1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 
    1014.57, 1014.59, 1014.61, 1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 
    1014.73, 1014.75, 1014.77, 1014.79, 1014.81, 1014.83,
  1014.3, 1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 
    1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 
    1014.62, 1014.64, 1014.66, 1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 
    1014.78, 1014.8, 1014.82, 1014.84, 1014.86, 1014.88,
  1014.35, 1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 
    1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 1014.63, 1014.65, 
    1014.67, 1014.69, 1014.71, 1014.73, 1014.75, 1014.77, 1014.79, 1014.81, 
    1014.83, 1014.85, 1014.87, 1014.89, 1014.91, 1014.93,
  1014.4, 1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 
    1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 1014.68, 1014.7, 
    1014.72, 1014.74, 1014.76, 1014.78, 1014.8, 1014.82, 1014.84, 1014.86, 
    1014.88, 1014.9, 1014.92, 1014.94, 1014.96, 1014.98,
  1013.55, 1013.57, 1013.59, 1013.61, 1013.63, 1013.65, 1013.67, 1013.69, 
    1013.71, 1013.73, 1013.75, 1013.77, 1013.79, 1013.81, 1013.83, 1013.85, 
    1013.87, 1013.89, 1013.91, 1013.93, 1013.95, 1013.97, 1013.99, 1014.01, 
    1014.03, 1014.05, 1014.07, 1014.09, 1014.11, 1014.13,
  1013.6, 1013.62, 1013.64, 1013.66, 1013.68, 1013.7, 1013.72, 1013.74, 
    1013.76, 1013.78, 1013.8, 1013.82, 1013.84, 1013.86, 1013.88, 1013.9, 
    1013.92, 1013.94, 1013.96, 1013.98, 1014, 1014.02, 1014.04, 1014.06, 
    1014.08, 1014.1, 1014.12, 1014.14, 1014.16, 1014.18,
  1013.65, 1013.67, 1013.69, 1013.71, 1013.73, 1013.75, 1013.77, 1013.79, 
    1013.81, 1013.83, 1013.85, 1013.87, 1013.89, 1013.91, 1013.93, 1013.95, 
    1013.97, 1013.99, 1014.01, 1014.03, 1014.05, 1014.07, 1014.09, 1014.11, 
    1014.13, 1014.15, 1014.17, 1014.19, 1014.21, 1014.23,
  1013.7, 1013.72, 1013.74, 1013.76, 1013.78, 1013.8, 1013.82, 1013.84, 
    1013.86, 1013.88, 1013.9, 1013.92, 1013.94, 1013.96, 1013.98, 1014, 
    1014.02, 1014.04, 1014.06, 1014.08, 1014.1, 1014.12, 1014.14, 1014.16, 
    1014.18, 1014.2, 1014.22, 1014.24, 1014.26, 1014.28,
  1013.75, 1013.77, 1013.79, 1013.81, 1013.83, 1013.85, 1013.87, 1013.89, 
    1013.91, 1013.93, 1013.95, 1013.97, 1013.99, 1014.01, 1014.03, 1014.05, 
    1014.07, 1014.09, 1014.11, 1014.13, 1014.15, 1014.17, 1014.19, 1014.21, 
    1014.23, 1014.25, 1014.27, 1014.29, 1014.31, 1014.33,
  1013.8, 1013.82, 1013.84, 1013.86, 1013.88, 1013.9, 1013.92, 1013.94, 
    1013.96, 1013.98, 1014, 1014.02, 1014.04, 1014.06, 1014.08, 1014.1, 
    1014.12, 1014.14, 1014.16, 1014.18, 1014.2, 1014.22, 1014.24, 1014.26, 
    1014.28, 1014.3, 1014.32, 1014.34, 1014.36, 1014.38,
  1013.85, 1013.87, 1013.89, 1013.91, 1013.93, 1013.95, 1013.97, 1013.99, 
    1014.01, 1014.03, 1014.05, 1014.07, 1014.09, 1014.11, 1014.13, 1014.15, 
    1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 1014.31, 
    1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 1014.43,
  1013.9, 1013.92, 1013.94, 1013.96, 1013.98, 1014, 1014.02, 1014.04, 
    1014.06, 1014.08, 1014.1, 1014.12, 1014.14, 1014.16, 1014.18, 1014.2, 
    1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 1014.36, 
    1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 1014.48,
  1013.95, 1013.97, 1013.99, 1014.01, 1014.03, 1014.05, 1014.07, 1014.09, 
    1014.11, 1014.13, 1014.15, 1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 
    1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 
    1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 1014.53,
  1014, 1014.02, 1014.04, 1014.06, 1014.08, 1014.1, 1014.12, 1014.14, 
    1014.16, 1014.18, 1014.2, 1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 
    1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 
    1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 1014.58,
  1014.05, 1014.07, 1014.09, 1014.11, 1014.13, 1014.15, 1014.17, 1014.19, 
    1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 
    1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 
    1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 1014.63,
  1014.1, 1014.12, 1014.14, 1014.16, 1014.18, 1014.2, 1014.22, 1014.24, 
    1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 
    1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 
    1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 1014.68,
  1014.15, 1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 
    1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 
    1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 
    1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 1014.73,
  1014.2, 1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 
    1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 
    1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 
    1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 1014.78,
  1014.25, 1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 
    1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 
    1014.57, 1014.59, 1014.61, 1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 
    1014.73, 1014.75, 1014.77, 1014.79, 1014.81, 1014.83,
  1014.3, 1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 
    1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 
    1014.62, 1014.64, 1014.66, 1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 
    1014.78, 1014.8, 1014.82, 1014.84, 1014.86, 1014.88,
  1014.35, 1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 
    1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 1014.63, 1014.65, 
    1014.67, 1014.69, 1014.71, 1014.73, 1014.75, 1014.77, 1014.79, 1014.81, 
    1014.83, 1014.85, 1014.87, 1014.89, 1014.91, 1014.93,
  1014.4, 1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 
    1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 1014.68, 1014.7, 
    1014.72, 1014.74, 1014.76, 1014.78, 1014.8, 1014.82, 1014.84, 1014.86, 
    1014.88, 1014.9, 1014.92, 1014.94, 1014.96, 1014.98,
  1014.45, 1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 
    1014.61, 1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 1014.73, 1014.75, 
    1014.77, 1014.79, 1014.81, 1014.83, 1014.85, 1014.87, 1014.89, 1014.91, 
    1014.93, 1014.95, 1014.97, 1014.99, 1015.01, 1015.03,
  1014.5, 1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 
    1014.66, 1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 1014.78, 1014.8, 
    1014.82, 1014.84, 1014.86, 1014.88, 1014.9, 1014.92, 1014.94, 1014.96, 
    1014.98, 1015, 1015.02, 1015.04, 1015.06, 1015.08,
  1013.65, 1013.67, 1013.69, 1013.71, 1013.73, 1013.75, 1013.77, 1013.79, 
    1013.81, 1013.83, 1013.85, 1013.87, 1013.89, 1013.91, 1013.93, 1013.95, 
    1013.97, 1013.99, 1014.01, 1014.03, 1014.05, 1014.07, 1014.09, 1014.11, 
    1014.13, 1014.15, 1014.17, 1014.19, 1014.21, 1014.23,
  1013.7, 1013.72, 1013.74, 1013.76, 1013.78, 1013.8, 1013.82, 1013.84, 
    1013.86, 1013.88, 1013.9, 1013.92, 1013.94, 1013.96, 1013.98, 1014, 
    1014.02, 1014.04, 1014.06, 1014.08, 1014.1, 1014.12, 1014.14, 1014.16, 
    1014.18, 1014.2, 1014.22, 1014.24, 1014.26, 1014.28,
  1013.75, 1013.77, 1013.79, 1013.81, 1013.83, 1013.85, 1013.87, 1013.89, 
    1013.91, 1013.93, 1013.95, 1013.97, 1013.99, 1014.01, 1014.03, 1014.05, 
    1014.07, 1014.09, 1014.11, 1014.13, 1014.15, 1014.17, 1014.19, 1014.21, 
    1014.23, 1014.25, 1014.27, 1014.29, 1014.31, 1014.33,
  1013.8, 1013.82, 1013.84, 1013.86, 1013.88, 1013.9, 1013.92, 1013.94, 
    1013.96, 1013.98, 1014, 1014.02, 1014.04, 1014.06, 1014.08, 1014.1, 
    1014.12, 1014.14, 1014.16, 1014.18, 1014.2, 1014.22, 1014.24, 1014.26, 
    1014.28, 1014.3, 1014.32, 1014.34, 1014.36, 1014.38,
  1013.85, 1013.87, 1013.89, 1013.91, 1013.93, 1013.95, 1013.97, 1013.99, 
    1014.01, 1014.03, 1014.05, 1014.07, 1014.09, 1014.11, 1014.13, 1014.15, 
    1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 1014.31, 
    1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 1014.43,
  1013.9, 1013.92, 1013.94, 1013.96, 1013.98, 1014, 1014.02, 1014.04, 
    1014.06, 1014.08, 1014.1, 1014.12, 1014.14, 1014.16, 1014.18, 1014.2, 
    1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 1014.36, 
    1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 1014.48,
  1013.95, 1013.97, 1013.99, 1014.01, 1014.03, 1014.05, 1014.07, 1014.09, 
    1014.11, 1014.13, 1014.15, 1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 
    1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 
    1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 1014.53,
  1014, 1014.02, 1014.04, 1014.06, 1014.08, 1014.1, 1014.12, 1014.14, 
    1014.16, 1014.18, 1014.2, 1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 
    1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 
    1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 1014.58,
  1014.05, 1014.07, 1014.09, 1014.11, 1014.13, 1014.15, 1014.17, 1014.19, 
    1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 
    1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 
    1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 1014.63,
  1014.1, 1014.12, 1014.14, 1014.16, 1014.18, 1014.2, 1014.22, 1014.24, 
    1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 
    1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 
    1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 1014.68,
  1014.15, 1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 
    1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 
    1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 
    1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 1014.73,
  1014.2, 1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 
    1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 
    1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 
    1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 1014.78,
  1014.25, 1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 
    1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 
    1014.57, 1014.59, 1014.61, 1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 
    1014.73, 1014.75, 1014.77, 1014.79, 1014.81, 1014.83,
  1014.3, 1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 
    1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 
    1014.62, 1014.64, 1014.66, 1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 
    1014.78, 1014.8, 1014.82, 1014.84, 1014.86, 1014.88,
  1014.35, 1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 
    1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 1014.63, 1014.65, 
    1014.67, 1014.69, 1014.71, 1014.73, 1014.75, 1014.77, 1014.79, 1014.81, 
    1014.83, 1014.85, 1014.87, 1014.89, 1014.91, 1014.93,
  1014.4, 1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 
    1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 1014.68, 1014.7, 
    1014.72, 1014.74, 1014.76, 1014.78, 1014.8, 1014.82, 1014.84, 1014.86, 
    1014.88, 1014.9, 1014.92, 1014.94, 1014.96, 1014.98,
  1014.45, 1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 
    1014.61, 1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 1014.73, 1014.75, 
    1014.77, 1014.79, 1014.81, 1014.83, 1014.85, 1014.87, 1014.89, 1014.91, 
    1014.93, 1014.95, 1014.97, 1014.99, 1015.01, 1015.03,
  1014.5, 1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 
    1014.66, 1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 1014.78, 1014.8, 
    1014.82, 1014.84, 1014.86, 1014.88, 1014.9, 1014.92, 1014.94, 1014.96, 
    1014.98, 1015, 1015.02, 1015.04, 1015.06, 1015.08,
  1014.55, 1014.57, 1014.59, 1014.61, 1014.63, 1014.65, 1014.67, 1014.69, 
    1014.71, 1014.73, 1014.75, 1014.77, 1014.79, 1014.81, 1014.83, 1014.85, 
    1014.87, 1014.89, 1014.91, 1014.93, 1014.95, 1014.97, 1014.99, 1015.01, 
    1015.03, 1015.05, 1015.07, 1015.09, 1015.11, 1015.13,
  1014.6, 1014.62, 1014.64, 1014.66, 1014.68, 1014.7, 1014.72, 1014.74, 
    1014.76, 1014.78, 1014.8, 1014.82, 1014.84, 1014.86, 1014.88, 1014.9, 
    1014.92, 1014.94, 1014.96, 1014.98, 1015, 1015.02, 1015.04, 1015.06, 
    1015.08, 1015.1, 1015.12, 1015.14, 1015.16, 1015.18,
  1013.75, 1013.77, 1013.79, 1013.81, 1013.83, 1013.85, 1013.87, 1013.89, 
    1013.91, 1013.93, 1013.95, 1013.97, 1013.99, 1014.01, 1014.03, 1014.05, 
    1014.07, 1014.09, 1014.11, 1014.13, 1014.15, 1014.17, 1014.19, 1014.21, 
    1014.23, 1014.25, 1014.27, 1014.29, 1014.31, 1014.33,
  1013.8, 1013.82, 1013.84, 1013.86, 1013.88, 1013.9, 1013.92, 1013.94, 
    1013.96, 1013.98, 1014, 1014.02, 1014.04, 1014.06, 1014.08, 1014.1, 
    1014.12, 1014.14, 1014.16, 1014.18, 1014.2, 1014.22, 1014.24, 1014.26, 
    1014.28, 1014.3, 1014.32, 1014.34, 1014.36, 1014.38,
  1013.85, 1013.87, 1013.89, 1013.91, 1013.93, 1013.95, 1013.97, 1013.99, 
    1014.01, 1014.03, 1014.05, 1014.07, 1014.09, 1014.11, 1014.13, 1014.15, 
    1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 1014.31, 
    1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 1014.43,
  1013.9, 1013.92, 1013.94, 1013.96, 1013.98, 1014, 1014.02, 1014.04, 
    1014.06, 1014.08, 1014.1, 1014.12, 1014.14, 1014.16, 1014.18, 1014.2, 
    1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 1014.36, 
    1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 1014.48,
  1013.95, 1013.97, 1013.99, 1014.01, 1014.03, 1014.05, 1014.07, 1014.09, 
    1014.11, 1014.13, 1014.15, 1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 
    1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 
    1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 1014.53,
  1014, 1014.02, 1014.04, 1014.06, 1014.08, 1014.1, 1014.12, 1014.14, 
    1014.16, 1014.18, 1014.2, 1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 
    1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 
    1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 1014.58,
  1014.05, 1014.07, 1014.09, 1014.11, 1014.13, 1014.15, 1014.17, 1014.19, 
    1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 
    1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 
    1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 1014.63,
  1014.1, 1014.12, 1014.14, 1014.16, 1014.18, 1014.2, 1014.22, 1014.24, 
    1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 
    1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 
    1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 1014.68,
  1014.15, 1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 
    1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 
    1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 
    1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 1014.73,
  1014.2, 1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 
    1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 
    1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 
    1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 1014.78,
  1014.25, 1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 
    1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 
    1014.57, 1014.59, 1014.61, 1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 
    1014.73, 1014.75, 1014.77, 1014.79, 1014.81, 1014.83,
  1014.3, 1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 
    1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 
    1014.62, 1014.64, 1014.66, 1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 
    1014.78, 1014.8, 1014.82, 1014.84, 1014.86, 1014.88,
  1014.35, 1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 
    1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 1014.63, 1014.65, 
    1014.67, 1014.69, 1014.71, 1014.73, 1014.75, 1014.77, 1014.79, 1014.81, 
    1014.83, 1014.85, 1014.87, 1014.89, 1014.91, 1014.93,
  1014.4, 1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 
    1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 1014.68, 1014.7, 
    1014.72, 1014.74, 1014.76, 1014.78, 1014.8, 1014.82, 1014.84, 1014.86, 
    1014.88, 1014.9, 1014.92, 1014.94, 1014.96, 1014.98,
  1014.45, 1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 
    1014.61, 1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 1014.73, 1014.75, 
    1014.77, 1014.79, 1014.81, 1014.83, 1014.85, 1014.87, 1014.89, 1014.91, 
    1014.93, 1014.95, 1014.97, 1014.99, 1015.01, 1015.03,
  1014.5, 1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 
    1014.66, 1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 1014.78, 1014.8, 
    1014.82, 1014.84, 1014.86, 1014.88, 1014.9, 1014.92, 1014.94, 1014.96, 
    1014.98, 1015, 1015.02, 1015.04, 1015.06, 1015.08,
  1014.55, 1014.57, 1014.59, 1014.61, 1014.63, 1014.65, 1014.67, 1014.69, 
    1014.71, 1014.73, 1014.75, 1014.77, 1014.79, 1014.81, 1014.83, 1014.85, 
    1014.87, 1014.89, 1014.91, 1014.93, 1014.95, 1014.97, 1014.99, 1015.01, 
    1015.03, 1015.05, 1015.07, 1015.09, 1015.11, 1015.13,
  1014.6, 1014.62, 1014.64, 1014.66, 1014.68, 1014.7, 1014.72, 1014.74, 
    1014.76, 1014.78, 1014.8, 1014.82, 1014.84, 1014.86, 1014.88, 1014.9, 
    1014.92, 1014.94, 1014.96, 1014.98, 1015, 1015.02, 1015.04, 1015.06, 
    1015.08, 1015.1, 1015.12, 1015.14, 1015.16, 1015.18,
  1014.65, 1014.67, 1014.69, 1014.71, 1014.73, 1014.75, 1014.77, 1014.79, 
    1014.81, 1014.83, 1014.85, 1014.87, 1014.89, 1014.91, 1014.93, 1014.95, 
    1014.97, 1014.99, 1015.01, 1015.03, 1015.05, 1015.07, 1015.09, 1015.11, 
    1015.13, 1015.15, 1015.17, 1015.19, 1015.21, 1015.23,
  1014.7, 1014.72, 1014.74, 1014.76, 1014.78, 1014.8, 1014.82, 1014.84, 
    1014.86, 1014.88, 1014.9, 1014.92, 1014.94, 1014.96, 1014.98, 1015, 
    1015.02, 1015.04, 1015.06, 1015.08, 1015.1, 1015.12, 1015.14, 1015.16, 
    1015.18, 1015.2, 1015.22, 1015.24, 1015.26, 1015.28,
  1013.85, 1013.87, 1013.89, 1013.91, 1013.93, 1013.95, 1013.97, 1013.99, 
    1014.01, 1014.03, 1014.05, 1014.07, 1014.09, 1014.11, 1014.13, 1014.15, 
    1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 1014.31, 
    1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 1014.43,
  1013.9, 1013.92, 1013.94, 1013.96, 1013.98, 1014, 1014.02, 1014.04, 
    1014.06, 1014.08, 1014.1, 1014.12, 1014.14, 1014.16, 1014.18, 1014.2, 
    1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 1014.36, 
    1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 1014.48,
  1013.95, 1013.97, 1013.99, 1014.01, 1014.03, 1014.05, 1014.07, 1014.09, 
    1014.11, 1014.13, 1014.15, 1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 
    1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 
    1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 1014.53,
  1014, 1014.02, 1014.04, 1014.06, 1014.08, 1014.1, 1014.12, 1014.14, 
    1014.16, 1014.18, 1014.2, 1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 
    1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 
    1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 1014.58,
  1014.05, 1014.07, 1014.09, 1014.11, 1014.13, 1014.15, 1014.17, 1014.19, 
    1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 
    1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 
    1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 1014.63,
  1014.1, 1014.12, 1014.14, 1014.16, 1014.18, 1014.2, 1014.22, 1014.24, 
    1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 
    1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 
    1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 1014.68,
  1014.15, 1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 
    1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 
    1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 
    1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 1014.73,
  1014.2, 1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 
    1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 
    1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 
    1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 1014.78,
  1014.25, 1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 
    1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 
    1014.57, 1014.59, 1014.61, 1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 
    1014.73, 1014.75, 1014.77, 1014.79, 1014.81, 1014.83,
  1014.3, 1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 
    1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 
    1014.62, 1014.64, 1014.66, 1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 
    1014.78, 1014.8, 1014.82, 1014.84, 1014.86, 1014.88,
  1014.35, 1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 
    1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 1014.63, 1014.65, 
    1014.67, 1014.69, 1014.71, 1014.73, 1014.75, 1014.77, 1014.79, 1014.81, 
    1014.83, 1014.85, 1014.87, 1014.89, 1014.91, 1014.93,
  1014.4, 1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 
    1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 1014.68, 1014.7, 
    1014.72, 1014.74, 1014.76, 1014.78, 1014.8, 1014.82, 1014.84, 1014.86, 
    1014.88, 1014.9, 1014.92, 1014.94, 1014.96, 1014.98,
  1014.45, 1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 
    1014.61, 1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 1014.73, 1014.75, 
    1014.77, 1014.79, 1014.81, 1014.83, 1014.85, 1014.87, 1014.89, 1014.91, 
    1014.93, 1014.95, 1014.97, 1014.99, 1015.01, 1015.03,
  1014.5, 1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 
    1014.66, 1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 1014.78, 1014.8, 
    1014.82, 1014.84, 1014.86, 1014.88, 1014.9, 1014.92, 1014.94, 1014.96, 
    1014.98, 1015, 1015.02, 1015.04, 1015.06, 1015.08,
  1014.55, 1014.57, 1014.59, 1014.61, 1014.63, 1014.65, 1014.67, 1014.69, 
    1014.71, 1014.73, 1014.75, 1014.77, 1014.79, 1014.81, 1014.83, 1014.85, 
    1014.87, 1014.89, 1014.91, 1014.93, 1014.95, 1014.97, 1014.99, 1015.01, 
    1015.03, 1015.05, 1015.07, 1015.09, 1015.11, 1015.13,
  1014.6, 1014.62, 1014.64, 1014.66, 1014.68, 1014.7, 1014.72, 1014.74, 
    1014.76, 1014.78, 1014.8, 1014.82, 1014.84, 1014.86, 1014.88, 1014.9, 
    1014.92, 1014.94, 1014.96, 1014.98, 1015, 1015.02, 1015.04, 1015.06, 
    1015.08, 1015.1, 1015.12, 1015.14, 1015.16, 1015.18,
  1014.65, 1014.67, 1014.69, 1014.71, 1014.73, 1014.75, 1014.77, 1014.79, 
    1014.81, 1014.83, 1014.85, 1014.87, 1014.89, 1014.91, 1014.93, 1014.95, 
    1014.97, 1014.99, 1015.01, 1015.03, 1015.05, 1015.07, 1015.09, 1015.11, 
    1015.13, 1015.15, 1015.17, 1015.19, 1015.21, 1015.23,
  1014.7, 1014.72, 1014.74, 1014.76, 1014.78, 1014.8, 1014.82, 1014.84, 
    1014.86, 1014.88, 1014.9, 1014.92, 1014.94, 1014.96, 1014.98, 1015, 
    1015.02, 1015.04, 1015.06, 1015.08, 1015.1, 1015.12, 1015.14, 1015.16, 
    1015.18, 1015.2, 1015.22, 1015.24, 1015.26, 1015.28,
  1014.75, 1014.77, 1014.79, 1014.81, 1014.83, 1014.85, 1014.87, 1014.89, 
    1014.91, 1014.93, 1014.95, 1014.97, 1014.99, 1015.01, 1015.03, 1015.05, 
    1015.07, 1015.09, 1015.11, 1015.13, 1015.15, 1015.17, 1015.19, 1015.21, 
    1015.23, 1015.25, 1015.27, 1015.29, 1015.31, 1015.33,
  1014.8, 1014.82, 1014.84, 1014.86, 1014.88, 1014.9, 1014.92, 1014.94, 
    1014.96, 1014.98, 1015, 1015.02, 1015.04, 1015.06, 1015.08, 1015.1, 
    1015.12, 1015.14, 1015.16, 1015.18, 1015.2, 1015.22, 1015.24, 1015.26, 
    1015.28, 1015.3, 1015.32, 1015.34, 1015.36, 1015.38,
  1013.95, 1013.97, 1013.99, 1014.01, 1014.03, 1014.05, 1014.07, 1014.09, 
    1014.11, 1014.13, 1014.15, 1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 
    1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 
    1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 1014.53,
  1014, 1014.02, 1014.04, 1014.06, 1014.08, 1014.1, 1014.12, 1014.14, 
    1014.16, 1014.18, 1014.2, 1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 
    1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 
    1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 1014.58,
  1014.05, 1014.07, 1014.09, 1014.11, 1014.13, 1014.15, 1014.17, 1014.19, 
    1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 
    1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 
    1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 1014.63,
  1014.1, 1014.12, 1014.14, 1014.16, 1014.18, 1014.2, 1014.22, 1014.24, 
    1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 
    1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 
    1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 1014.68,
  1014.15, 1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 
    1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 
    1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 
    1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 1014.73,
  1014.2, 1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 
    1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 
    1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 
    1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 1014.78,
  1014.25, 1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 
    1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 
    1014.57, 1014.59, 1014.61, 1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 
    1014.73, 1014.75, 1014.77, 1014.79, 1014.81, 1014.83,
  1014.3, 1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 
    1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 
    1014.62, 1014.64, 1014.66, 1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 
    1014.78, 1014.8, 1014.82, 1014.84, 1014.86, 1014.88,
  1014.35, 1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 
    1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 1014.63, 1014.65, 
    1014.67, 1014.69, 1014.71, 1014.73, 1014.75, 1014.77, 1014.79, 1014.81, 
    1014.83, 1014.85, 1014.87, 1014.89, 1014.91, 1014.93,
  1014.4, 1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 
    1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 1014.68, 1014.7, 
    1014.72, 1014.74, 1014.76, 1014.78, 1014.8, 1014.82, 1014.84, 1014.86, 
    1014.88, 1014.9, 1014.92, 1014.94, 1014.96, 1014.98,
  1014.45, 1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 
    1014.61, 1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 1014.73, 1014.75, 
    1014.77, 1014.79, 1014.81, 1014.83, 1014.85, 1014.87, 1014.89, 1014.91, 
    1014.93, 1014.95, 1014.97, 1014.99, 1015.01, 1015.03,
  1014.5, 1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 
    1014.66, 1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 1014.78, 1014.8, 
    1014.82, 1014.84, 1014.86, 1014.88, 1014.9, 1014.92, 1014.94, 1014.96, 
    1014.98, 1015, 1015.02, 1015.04, 1015.06, 1015.08,
  1014.55, 1014.57, 1014.59, 1014.61, 1014.63, 1014.65, 1014.67, 1014.69, 
    1014.71, 1014.73, 1014.75, 1014.77, 1014.79, 1014.81, 1014.83, 1014.85, 
    1014.87, 1014.89, 1014.91, 1014.93, 1014.95, 1014.97, 1014.99, 1015.01, 
    1015.03, 1015.05, 1015.07, 1015.09, 1015.11, 1015.13,
  1014.6, 1014.62, 1014.64, 1014.66, 1014.68, 1014.7, 1014.72, 1014.74, 
    1014.76, 1014.78, 1014.8, 1014.82, 1014.84, 1014.86, 1014.88, 1014.9, 
    1014.92, 1014.94, 1014.96, 1014.98, 1015, 1015.02, 1015.04, 1015.06, 
    1015.08, 1015.1, 1015.12, 1015.14, 1015.16, 1015.18,
  1014.65, 1014.67, 1014.69, 1014.71, 1014.73, 1014.75, 1014.77, 1014.79, 
    1014.81, 1014.83, 1014.85, 1014.87, 1014.89, 1014.91, 1014.93, 1014.95, 
    1014.97, 1014.99, 1015.01, 1015.03, 1015.05, 1015.07, 1015.09, 1015.11, 
    1015.13, 1015.15, 1015.17, 1015.19, 1015.21, 1015.23,
  1014.7, 1014.72, 1014.74, 1014.76, 1014.78, 1014.8, 1014.82, 1014.84, 
    1014.86, 1014.88, 1014.9, 1014.92, 1014.94, 1014.96, 1014.98, 1015, 
    1015.02, 1015.04, 1015.06, 1015.08, 1015.1, 1015.12, 1015.14, 1015.16, 
    1015.18, 1015.2, 1015.22, 1015.24, 1015.26, 1015.28,
  1014.75, 1014.77, 1014.79, 1014.81, 1014.83, 1014.85, 1014.87, 1014.89, 
    1014.91, 1014.93, 1014.95, 1014.97, 1014.99, 1015.01, 1015.03, 1015.05, 
    1015.07, 1015.09, 1015.11, 1015.13, 1015.15, 1015.17, 1015.19, 1015.21, 
    1015.23, 1015.25, 1015.27, 1015.29, 1015.31, 1015.33,
  1014.8, 1014.82, 1014.84, 1014.86, 1014.88, 1014.9, 1014.92, 1014.94, 
    1014.96, 1014.98, 1015, 1015.02, 1015.04, 1015.06, 1015.08, 1015.1, 
    1015.12, 1015.14, 1015.16, 1015.18, 1015.2, 1015.22, 1015.24, 1015.26, 
    1015.28, 1015.3, 1015.32, 1015.34, 1015.36, 1015.38,
  1014.85, 1014.87, 1014.89, 1014.91, 1014.93, 1014.95, 1014.97, 1014.99, 
    1015.01, 1015.03, 1015.05, 1015.07, 1015.09, 1015.11, 1015.13, 1015.15, 
    1015.17, 1015.19, 1015.21, 1015.23, 1015.25, 1015.27, 1015.29, 1015.31, 
    1015.33, 1015.35, 1015.37, 1015.39, 1015.41, 1015.43,
  1014.9, 1014.92, 1014.94, 1014.96, 1014.98, 1015, 1015.02, 1015.04, 
    1015.06, 1015.08, 1015.1, 1015.12, 1015.14, 1015.16, 1015.18, 1015.2, 
    1015.22, 1015.24, 1015.26, 1015.28, 1015.3, 1015.32, 1015.34, 1015.36, 
    1015.38, 1015.4, 1015.42, 1015.44, 1015.46, 1015.48,
  1014.05, 1014.07, 1014.09, 1014.11, 1014.13, 1014.15, 1014.17, 1014.19, 
    1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 
    1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 
    1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 1014.63,
  1014.1, 1014.12, 1014.14, 1014.16, 1014.18, 1014.2, 1014.22, 1014.24, 
    1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 
    1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 
    1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 1014.68,
  1014.15, 1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 
    1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 
    1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 
    1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 1014.73,
  1014.2, 1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 
    1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 
    1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 
    1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 1014.78,
  1014.25, 1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 
    1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 
    1014.57, 1014.59, 1014.61, 1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 
    1014.73, 1014.75, 1014.77, 1014.79, 1014.81, 1014.83,
  1014.3, 1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 
    1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 
    1014.62, 1014.64, 1014.66, 1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 
    1014.78, 1014.8, 1014.82, 1014.84, 1014.86, 1014.88,
  1014.35, 1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 
    1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 1014.63, 1014.65, 
    1014.67, 1014.69, 1014.71, 1014.73, 1014.75, 1014.77, 1014.79, 1014.81, 
    1014.83, 1014.85, 1014.87, 1014.89, 1014.91, 1014.93,
  1014.4, 1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 
    1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 1014.68, 1014.7, 
    1014.72, 1014.74, 1014.76, 1014.78, 1014.8, 1014.82, 1014.84, 1014.86, 
    1014.88, 1014.9, 1014.92, 1014.94, 1014.96, 1014.98,
  1014.45, 1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 
    1014.61, 1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 1014.73, 1014.75, 
    1014.77, 1014.79, 1014.81, 1014.83, 1014.85, 1014.87, 1014.89, 1014.91, 
    1014.93, 1014.95, 1014.97, 1014.99, 1015.01, 1015.03,
  1014.5, 1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 
    1014.66, 1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 1014.78, 1014.8, 
    1014.82, 1014.84, 1014.86, 1014.88, 1014.9, 1014.92, 1014.94, 1014.96, 
    1014.98, 1015, 1015.02, 1015.04, 1015.06, 1015.08,
  1014.55, 1014.57, 1014.59, 1014.61, 1014.63, 1014.65, 1014.67, 1014.69, 
    1014.71, 1014.73, 1014.75, 1014.77, 1014.79, 1014.81, 1014.83, 1014.85, 
    1014.87, 1014.89, 1014.91, 1014.93, 1014.95, 1014.97, 1014.99, 1015.01, 
    1015.03, 1015.05, 1015.07, 1015.09, 1015.11, 1015.13,
  1014.6, 1014.62, 1014.64, 1014.66, 1014.68, 1014.7, 1014.72, 1014.74, 
    1014.76, 1014.78, 1014.8, 1014.82, 1014.84, 1014.86, 1014.88, 1014.9, 
    1014.92, 1014.94, 1014.96, 1014.98, 1015, 1015.02, 1015.04, 1015.06, 
    1015.08, 1015.1, 1015.12, 1015.14, 1015.16, 1015.18,
  1014.65, 1014.67, 1014.69, 1014.71, 1014.73, 1014.75, 1014.77, 1014.79, 
    1014.81, 1014.83, 1014.85, 1014.87, 1014.89, 1014.91, 1014.93, 1014.95, 
    1014.97, 1014.99, 1015.01, 1015.03, 1015.05, 1015.07, 1015.09, 1015.11, 
    1015.13, 1015.15, 1015.17, 1015.19, 1015.21, 1015.23,
  1014.7, 1014.72, 1014.74, 1014.76, 1014.78, 1014.8, 1014.82, 1014.84, 
    1014.86, 1014.88, 1014.9, 1014.92, 1014.94, 1014.96, 1014.98, 1015, 
    1015.02, 1015.04, 1015.06, 1015.08, 1015.1, 1015.12, 1015.14, 1015.16, 
    1015.18, 1015.2, 1015.22, 1015.24, 1015.26, 1015.28,
  1014.75, 1014.77, 1014.79, 1014.81, 1014.83, 1014.85, 1014.87, 1014.89, 
    1014.91, 1014.93, 1014.95, 1014.97, 1014.99, 1015.01, 1015.03, 1015.05, 
    1015.07, 1015.09, 1015.11, 1015.13, 1015.15, 1015.17, 1015.19, 1015.21, 
    1015.23, 1015.25, 1015.27, 1015.29, 1015.31, 1015.33,
  1014.8, 1014.82, 1014.84, 1014.86, 1014.88, 1014.9, 1014.92, 1014.94, 
    1014.96, 1014.98, 1015, 1015.02, 1015.04, 1015.06, 1015.08, 1015.1, 
    1015.12, 1015.14, 1015.16, 1015.18, 1015.2, 1015.22, 1015.24, 1015.26, 
    1015.28, 1015.3, 1015.32, 1015.34, 1015.36, 1015.38,
  1014.85, 1014.87, 1014.89, 1014.91, 1014.93, 1014.95, 1014.97, 1014.99, 
    1015.01, 1015.03, 1015.05, 1015.07, 1015.09, 1015.11, 1015.13, 1015.15, 
    1015.17, 1015.19, 1015.21, 1015.23, 1015.25, 1015.27, 1015.29, 1015.31, 
    1015.33, 1015.35, 1015.37, 1015.39, 1015.41, 1015.43,
  1014.9, 1014.92, 1014.94, 1014.96, 1014.98, 1015, 1015.02, 1015.04, 
    1015.06, 1015.08, 1015.1, 1015.12, 1015.14, 1015.16, 1015.18, 1015.2, 
    1015.22, 1015.24, 1015.26, 1015.28, 1015.3, 1015.32, 1015.34, 1015.36, 
    1015.38, 1015.4, 1015.42, 1015.44, 1015.46, 1015.48,
  1014.95, 1014.97, 1014.99, 1015.01, 1015.03, 1015.05, 1015.07, 1015.09, 
    1015.11, 1015.13, 1015.15, 1015.17, 1015.19, 1015.21, 1015.23, 1015.25, 
    1015.27, 1015.29, 1015.31, 1015.33, 1015.35, 1015.37, 1015.39, 1015.41, 
    1015.43, 1015.45, 1015.47, 1015.49, 1015.51, 1015.53,
  1015, 1015.02, 1015.04, 1015.06, 1015.08, 1015.1, 1015.12, 1015.14, 
    1015.16, 1015.18, 1015.2, 1015.22, 1015.24, 1015.26, 1015.28, 1015.3, 
    1015.32, 1015.34, 1015.36, 1015.38, 1015.4, 1015.42, 1015.44, 1015.46, 
    1015.48, 1015.5, 1015.52, 1015.54, 1015.56, 1015.58,
  1014.15, 1014.17, 1014.19, 1014.21, 1014.23, 1014.25, 1014.27, 1014.29, 
    1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 
    1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 
    1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 1014.73,
  1014.2, 1014.22, 1014.24, 1014.26, 1014.28, 1014.3, 1014.32, 1014.34, 
    1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 
    1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 
    1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 1014.78,
  1014.25, 1014.27, 1014.29, 1014.31, 1014.33, 1014.35, 1014.37, 1014.39, 
    1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 
    1014.57, 1014.59, 1014.61, 1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 
    1014.73, 1014.75, 1014.77, 1014.79, 1014.81, 1014.83,
  1014.3, 1014.32, 1014.34, 1014.36, 1014.38, 1014.4, 1014.42, 1014.44, 
    1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 
    1014.62, 1014.64, 1014.66, 1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 
    1014.78, 1014.8, 1014.82, 1014.84, 1014.86, 1014.88,
  1014.35, 1014.37, 1014.39, 1014.41, 1014.43, 1014.45, 1014.47, 1014.49, 
    1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 1014.61, 1014.63, 1014.65, 
    1014.67, 1014.69, 1014.71, 1014.73, 1014.75, 1014.77, 1014.79, 1014.81, 
    1014.83, 1014.85, 1014.87, 1014.89, 1014.91, 1014.93,
  1014.4, 1014.42, 1014.44, 1014.46, 1014.48, 1014.5, 1014.52, 1014.54, 
    1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 1014.66, 1014.68, 1014.7, 
    1014.72, 1014.74, 1014.76, 1014.78, 1014.8, 1014.82, 1014.84, 1014.86, 
    1014.88, 1014.9, 1014.92, 1014.94, 1014.96, 1014.98,
  1014.45, 1014.47, 1014.49, 1014.51, 1014.53, 1014.55, 1014.57, 1014.59, 
    1014.61, 1014.63, 1014.65, 1014.67, 1014.69, 1014.71, 1014.73, 1014.75, 
    1014.77, 1014.79, 1014.81, 1014.83, 1014.85, 1014.87, 1014.89, 1014.91, 
    1014.93, 1014.95, 1014.97, 1014.99, 1015.01, 1015.03,
  1014.5, 1014.52, 1014.54, 1014.56, 1014.58, 1014.6, 1014.62, 1014.64, 
    1014.66, 1014.68, 1014.7, 1014.72, 1014.74, 1014.76, 1014.78, 1014.8, 
    1014.82, 1014.84, 1014.86, 1014.88, 1014.9, 1014.92, 1014.94, 1014.96, 
    1014.98, 1015, 1015.02, 1015.04, 1015.06, 1015.08,
  1014.55, 1014.57, 1014.59, 1014.61, 1014.63, 1014.65, 1014.67, 1014.69, 
    1014.71, 1014.73, 1014.75, 1014.77, 1014.79, 1014.81, 1014.83, 1014.85, 
    1014.87, 1014.89, 1014.91, 1014.93, 1014.95, 1014.97, 1014.99, 1015.01, 
    1015.03, 1015.05, 1015.07, 1015.09, 1015.11, 1015.13,
  1014.6, 1014.62, 1014.64, 1014.66, 1014.68, 1014.7, 1014.72, 1014.74, 
    1014.76, 1014.78, 1014.8, 1014.82, 1014.84, 1014.86, 1014.88, 1014.9, 
    1014.92, 1014.94, 1014.96, 1014.98, 1015, 1015.02, 1015.04, 1015.06, 
    1015.08, 1015.1, 1015.12, 1015.14, 1015.16, 1015.18,
  1014.65, 1014.67, 1014.69, 1014.71, 1014.73, 1014.75, 1014.77, 1014.79, 
    1014.81, 1014.83, 1014.85, 1014.87, 1014.89, 1014.91, 1014.93, 1014.95, 
    1014.97, 1014.99, 1015.01, 1015.03, 1015.05, 1015.07, 1015.09, 1015.11, 
    1015.13, 1015.15, 1015.17, 1015.19, 1015.21, 1015.23,
  1014.7, 1014.72, 1014.74, 1014.76, 1014.78, 1014.8, 1014.82, 1014.84, 
    1014.86, 1014.88, 1014.9, 1014.92, 1014.94, 1014.96, 1014.98, 1015, 
    1015.02, 1015.04, 1015.06, 1015.08, 1015.1, 1015.12, 1015.14, 1015.16, 
    1015.18, 1015.2, 1015.22, 1015.24, 1015.26, 1015.28,
  1014.75, 1014.77, 1014.79, 1014.81, 1014.83, 1014.85, 1014.87, 1014.89, 
    1014.91, 1014.93, 1014.95, 1014.97, 1014.99, 1015.01, 1015.03, 1015.05, 
    1015.07, 1015.09, 1015.11, 1015.13, 1015.15, 1015.17, 1015.19, 1015.21, 
    1015.23, 1015.25, 1015.27, 1015.29, 1015.31, 1015.33,
  1014.8, 1014.82, 1014.84, 1014.86, 1014.88, 1014.9, 1014.92, 1014.94, 
    1014.96, 1014.98, 1015, 1015.02, 1015.04, 1015.06, 1015.08, 1015.1, 
    1015.12, 1015.14, 1015.16, 1015.18, 1015.2, 1015.22, 1015.24, 1015.26, 
    1015.28, 1015.3, 1015.32, 1015.34, 1015.36, 1015.38,
  1014.85, 1014.87, 1014.89, 1014.91, 1014.93, 1014.95, 1014.97, 1014.99, 
    1015.01, 1015.03, 1015.05, 1015.07, 1015.09, 1015.11, 1015.13, 1015.15, 
    1015.17, 1015.19, 1015.21, 1015.23, 1015.25, 1015.27, 1015.29, 1015.31, 
    1015.33, 1015.35, 1015.37, 1015.39, 1015.41, 1015.43,
  1014.9, 1014.92, 1014.94, 1014.96, 1014.98, 1015, 1015.02, 1015.04, 
    1015.06, 1015.08, 1015.1, 1015.12, 1015.14, 1015.16, 1015.18, 1015.2, 
    1015.22, 1015.24, 1015.26, 1015.28, 1015.3, 1015.32, 1015.34, 1015.36, 
    1015.38, 1015.4, 1015.42, 1015.44, 1015.46, 1015.48,
  1014.95, 1014.97, 1014.99, 1015.01, 1015.03, 1015.05, 1015.07, 1015.09, 
    1015.11, 1015.13, 1015.15, 1015.17, 1015.19, 1015.21, 1015.23, 1015.25, 
    1015.27, 1015.29, 1015.31, 1015.33, 1015.35, 1015.37, 1015.39, 1015.41, 
    1015.43, 1015.45, 1015.47, 1015.49, 1015.51, 1015.53,
  1015, 1015.02, 1015.04, 1015.06, 1015.08, 1015.1, 1015.12, 1015.14, 
    1015.16, 1015.18, 1015.2, 1015.22, 1015.24, 1015.26, 1015.28, 1015.3, 
    1015.32, 1015.34, 1015.36, 1015.38, 1015.4, 1015.42, 1015.44, 1015.46, 
    1015.48, 1015.5, 1015.52, 1015.54, 1015.56, 1015.58,
  1015.05, 1015.07, 1015.09, 1015.11, 1015.13, 1015.15, 1015.17, 1015.19, 
    1015.21, 1015.23, 1015.25, 1015.27, 1015.29, 1015.31, 1015.33, 1015.35, 
    1015.37, 1015.39, 1015.41, 1015.43, 1015.45, 1015.47, 1015.49, 1015.51, 
    1015.53, 1015.55, 1015.57, 1015.59, 1015.61, 1015.63,
  1015.1, 1015.12, 1015.14, 1015.16, 1015.18, 1015.2, 1015.22, 1015.24, 
    1015.26, 1015.28, 1015.3, 1015.32, 1015.34, 1015.36, 1015.38, 1015.4, 
    1015.42, 1015.44, 1015.46, 1015.48, 1015.5, 1015.52, 1015.54, 1015.56, 
    1015.58, 1015.6, 1015.62, 1015.64, 1015.66, 1015.68 ;
}
