netcdf f_user_types {
types:
  opaque(16) calibration_t ;
}
