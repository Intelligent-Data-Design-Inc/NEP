netcdf unlimited_dim {
dimensions:
	time = UNLIMITED ; // (5 currently)
	lat = 4 ;
	lon = 5 ;
variables:
	float time(time) ;
	float temperature(time, lat, lon) ;
data:

 time = 0, 1, 2, 3, 4 ;

 temperature =
  273.15, 275.15, 277.15, 279.15, 281.15,
  278.15, 280.15, 282.15, 284.15, 286.15,
  283.15, 285.15, 287.15, 289.15, 291.15,
  288.15, 290.15, 292.15, 294.15, 296.15,
  274.15, 276.15, 278.15, 280.15, 282.15,
  279.15, 281.15, 283.15, 285.15, 287.15,
  284.15, 286.15, 288.15, 290.15, 292.15,
  289.15, 291.15, 293.15, 295.15, 297.15,
  275.15, 277.15, 279.15, 281.15, 283.15,
  280.15, 282.15, 284.15, 286.15, 288.15,
  285.15, 287.15, 289.15, 291.15, 293.15,
  290.15, 292.15, 294.15, 296.15, 298.15,
  276.15, 278.15, 280.15, 282.15, 284.15,
  281.15, 283.15, 285.15, 287.15, 289.15,
  286.15, 288.15, 290.15, 292.15, 294.15,
  291.15, 293.15, 295.15, 297.15, 299.15,
  277.15, 279.15, 281.15, 283.15, 285.15,
  282.15, 284.15, 286.15, 288.15, 290.15,
  287.15, 289.15, 291.15, 293.15, 295.15,
  292.15, 294.15, 296.15, 298.15, 300.15 ;
}
