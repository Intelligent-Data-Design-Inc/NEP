netcdf user_types {
types:
  compound weather_obs_t {
    double time ;
    float temperature ;
    float pressure ;
    float humidity ;
  }; // weather_obs_t
  int(*) obs_per_day_t ;
  int enum cloud_cover_t {CLEAR = 0, PARTLY_CLOUDY = 1, CLOUDY = 2, 
      OVERCAST = 3} ;
  opaque(16) calibration_t ;
dimensions:
	obs = 5 ;
	day = 3 ;
variables:
	weather_obs_t observations(obs) ;
	obs_per_day_t obs_per_day(day) ;
	cloud_cover_t cloud_cover(obs) ;
	calibration_t calibration ;
data:

 observations = {1000, 20, 1013, 60}, {4600, 22, 1013.5, 55}, 
    {8200, 24, 1014, 50}, {11800, 26, 1014.5, 45}, {15400, 28, 1015, 40} ;

 obs_per_day = {10, 15, 20}, {12, 18, 22, 25}, {8, 14} ;

 cloud_cover = CLEAR, PARTLY_CLOUDY, CLOUDY, PARTLY_CLOUDY, OVERCAST ;

 calibration = 0X00112233445566778899AABBCCDDEEFF ;
}
