netcdf f_multi_unlimited {
dimensions:
	station = UNLIMITED ; // (5 currently)
	time = UNLIMITED ; // (8 currently)
variables:
	float temperature(station, time) ;
data:

 temperature =
  {20, 20.5, 21, 21.5, 22, 22.5, 23, 23.5},
  {22, 22.5, 23, 23.5, 24, 24.5, 25, 25.5},
  {24, 24.5, 25, 25.5, 26, 26.5, 27, 27.5},
  {26, 26.5, 27, 27.5, 28, 28.5, 29, 29.5},
  {28, 28.5, 29, 29.5, 30, 30.5, 31, 31.5} ;
}
